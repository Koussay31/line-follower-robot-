PK   �|�X�`���
  �q     cirkitFile.json�]�۸��J��2�K�r�d�@�]$h��"�De���SY�G������K<�s&؋��%�}%R��w��%���YU�έ>�n�n7�S�ɍ���|o�H��ͪ߮�w��&y�%l���c���n�q�~em����J!��u��BKfs]N��r�&O߾[�a9��N.'���VkV�M�T�4˥p,�R�ei�T������cɧ��O��	.��-�)�jҒ��,����4%�f��O�$�;H>=v�W�(kɚ�vL�2�r'�T��VB4s̃��cɧ��O�]�Te9ϙ��3UJǊ�4��mx*��s̃��cɧ��#Ǯpr��g8���s��@b���G�Ǒ�q$z|��\YZ��U&��ba2Vԩc�lx�i������ ��Jg�FW�zQ��u�e�,K��>M����zn���g��0ª\���R��W��b��E%KW����x9��3�A�3�A�3�A�3"��x�LŃ�g*D>S�@�`�Cr7W�@z$ys��f�ԍ�m�?�F��QHV4�cZ�*�rm��3w=H>=� �����s�OO=H����$���A��$���a�`�Cr7s���H�f�z��G�Ǒ�q$~ɟ@�'�uɟ@�'��	$ɟ@�'�������x�ڮ�2^L��?	*e$p$.2��	\��"	\���%	\��)	\���,	\��0	\���3	\��7	\h�E��h���Ő��$.uD����i��4�r�y�`h|J�_��a*�K�`�J�Bs.q|�y+�K^`�J����,��%^}��,uD������Ԗ�x��F�.��v	\�W	���\�h��f�.�*M�)�#����x���64 UN�0�a��@�i(4�LC���X�P,h(4����S8��m������ή��4�E��Ș8�ƻD�N�]����.�y��x�輀�i�Kt^��4�%:/�p��p8�w��E�I\2C⒓�4��KC/������i �Q���4�%�ZC�i�K�h8�w�9�8��p��N�]��N�]��NPG/����	lh �W_p8�w�^'p8�w�^%p8�w��F�*��.�*�	�#����x����64 UN�0�a��@�i(4�LC���X�P,h(4������S�����?��c۹��n�?gիv��v��_�>4u�v����M}����}�9F���m�$�<|���4|���1z���i=8���g�N�1����m�~f��D��?8���g�N�1����j�~f����ǎ_!��ϐz���H}�� �@�E�c�X���4��[�	2F?� 45��ǟC�c�s Bsa�~�
B�`�~�
B�_?h ��VAp΋2�B8W��.F?s�I.F?s��-F����* �j1��* �gQ���8W�9,� !�
p,��!ǂȱ$
,�]�$
,�K���(�$
,�K�8��u���mrK��%$�K��M�W��	���;��]Br��BH sU��P�H�i�����W�_E�3t=y��C_:�����v:\�J�g��y�p@Ԩ����П
b�
"(DP��A!��C���� �������7Vƽ}���ږn��n�^���ٺ��.�"�ٮ��?�&`��x[�~������^u�;����ۻM�'���v��]�y��sco�vh]$�z�^��u���_t�ē_~~����-��v7ۏ/7�����]�oܹ�M�k˵;����m�<}�w~t�v������usgr��tJ����'Ϗ�$8��lwm?�Y�2K#
�P�M(8~Z�	��ݓ<׎g�a�q���`�;�d��]SE��]�7ǿ�H|���:���"�v�w��SK�w���/��,K���&���~�m��A�{ۿ��u�=�]r)}]�����K*�.���7',�\t~�?����c����.�g .ڜ������:ۯ~T��Å��z���"Ϊ���2=��|�*N����=:L<�~�Vۦ۷���z4� |��I����J��>̴:'���*OT�]�L�kL�YiK��<5bx��� �3�?�Q~��1���ЩHs9�6��G��M�L6bt���I��y"Z9�Փg��iU>�*��Ʉz3�$&�8,��zB�G��K�Y�c��Y��K�/�N��n���9�U�U&���ٰLˌ�BXfL#����,@��>Wg��K��U�Z��)��~E1�}�u1�P���Й�(SJ�Oa���y8�j�}&n�P���8����?^>c\���'X[^�������%�%��s�`���Ŋ�s�?Ц�Ii
�s�����FjYf���L�VH����-�{g}(�pX]�z��G�i�C𨇌z�k���m��<�]=�����ksuNƶ�3:�=��Q�b)��l��4�Z��U^�%��Ovμ/j�H+�ٴ���.kVX��-��2��'ƙ������������߹�Q��E�X��\;��r��J���bGxl(&N@�G~����W�ؘg�s�N�Ҝ?j�;i~��_T�m�>�����u�vh:��a˜�(}�vu؇&��U�x��l��V������ez�1\��-}:a����^�l)/a��;!���7��F�[��$L�49�ª�vMXsX���$|ս�o���ťV�;o\��&t婑�<|��t_��� �H��q��c��s}��M�>�+|�~����e��]���͛|�-��]��_;�����E�nw���?�]������ܮ�ڻ��J��PK   �|�XG�~��  � /   images/0739a1b1-a163-452a-a325-ab452d55b136.png�y8�m?�r�J�M!*IY��Ie�^Y&������[�d�cb�0��d�1̒,�ٲ�L������������|�|�4}��>�r}��|��mn$�_l��mۄ�o^�ܶM�i۶]&{w-�����A���{����� ��n�m�&�I����em4�6�l����
�*y�����x(����WŶm;����5��9t4Gb&��Ȳѹ�}��OܜΉSٱ������b��MT�}�L�1HƸD���?j��i͘�ǰf�	�A��{�ξ�[_����J�z���r���٢w��/5a��t�I��ե�EnhǶ-?����'m�ں-��Ǔ[�n�-��v<����xN��J�h���e3��2������7��=V��)u!";G?�� ��<�|K0�yY���I2,���^)�Ϭ���Ev�p�����������d���4���dK;!-�L�^�$Cx�䐦W��k��E���9謗	* P��ϕ�����S�����0C���~�?��$Ǖ���φ%mXJ����{���w/�y|
�T!��;��G����쳄�[�����⩧�U�6}3���6��{�[$��ab1�P��~z�3������Y�q(�V�f��¦�&	�� ��l.Z��s9�2SH�W�ơP6�[��SnT�QokF!s�Ǔ`��� 6rl�������fI�:�v�K�|l��%����)�m����}gw0�6=y�dk��?�/������<�w�}l��جJ���s�+����������6����Í�͍{3�����"R-33�	a\yoU+����̡-�߶~�S���v�ѯ�f��nY7�߼�K�pE߬�����f�J�\t���+"D�,�����AGf�H��X��i���&���oց���A{10�^���l����UL&0���ٵ?���E�)�Q�5��s�=[�,�8�v�Y����>\��>\+sS�N��88y��</�!-Ot�HS�/'9��q�ZwuR��
���ӝ�v�����xS>edf5�Ի`��Z��/�j�3�QM�/
�1Q �wH����G�h�p���"[�|���fi�h.��-
��f�:�[<?>gh8)�2d����q���j�GZl��Ϩ�4.{��F���Hq���5�1͸�m2�2~�l����]I���J�&k�-�x�T�/�O�z�5�k����8��JdX��a9�<��V��\�����R��9�����0�TƦ%r�hm�[o���b�Pԓ��YپQ5Y�� �>[Զ�f�UG~����bhA�A	���6��,-��:[��Y����p���m���k���A��p�ʂ�K��&�{sdJ;?=3�O�	}�Ij�>>wE�Ws20NJ]=X�uq�g�j����bN���|�G����Q�s˪�r���W��ӕ������7�[����v�ЂF�K^��FY�{��s��ʻ��R�:i��D{��x�����T�Dr��j�M�s3�����:u˙��[�.�[Im}�v8��0��d�Y�S�ܷ�BW�V�F��V�E��V�
���355;����҈�RW&/�+�'��]W�e����v�@$�Y��=�Vܲܽ��ٳ�6�tinb��[s!ޞ�C����<_��iG�Gn���_a+*�� ]>��-u��{\lrǹ��x�|�b�ߕ��?e��@�㕸�����[�`J�p-��i��m�'���n��:l�xm�pd�l�em,W0Q�:��"�A�fXDyP��pOTG^uPiN��c��+l����~ŭdyώ�ȂrZ�����?���A�Xc|O���/�Pc���>���tx/��g�N8^xai=���
\�ΟNXi��@�l��]Q�0��!a�+ץ���q�����`Vq,�o"�B8a�i���Itq�����1C�06�J��J���
�<-VTy�����kQ
�ɍ������p�F����Ϝ����r�}��O��u�~�Ar�u�����Wc~2�ƪ����@�m�����
&�H�;7��.2g�>)l!�(�|�v�z��[�TJ�й��#�J�:F���R���:oȼ�>33�w��vå"����P|�?{�&��#�H��+���#��<o��Jڐ(-�������&�Mt^��R��|٢����q`�g��c��j��02���)����F�;W������+�xR��:P��/�ސc�H���\k�Ý�/���d�����^� u �Ƚ���c��������-6yK�.�d�j��܉�x�������7�.{��"�'�>����K�۰o�g����m%���UY�> �/��
zo��X{_�v��Kû��q��Ŧ�ү2#G�_Z&�k3��x��r��2#zל���@�[��װ��^_�L�#/=lql�X4Xm������nq�p�7ME]�A��J60��e��ogU.Ė�FՄ�W_Ћ�[cT���l�hze< &��x����/{�"�Lv��
��= з$:��Ln�_�|_�!��ɬK{U���G��Jak�6����������R3Ć��S�ۿE$��|��ӝ1��E}��q[s<w�R��.�$����V�P���Lկ�0e�YK�9��qO_L���p��Tu��/8�ˊ��Z��]��A�@(�^�1���s�z��'�l��x�}u��A���<�� m������j��1õ��B��iB��	�A&q��6�t���+�cQ"M	��յN�I/&�'9�˹��Vv�t�R��FAD�/��"������N��+�',��Z.����xT�;(a��C��?����Drɴ��J@a��m�e��h?-����b	���M8=�^����=�ӽ�b/��Y:#�3���rp`��$G7��0_��s�N���vo���B��
]\�R�	�e�1cٝ)z)A���۹����E;DO�V$���t+˾C��@;�sA����.���8yQ\��Gwz�O/9s>u��ř����e�5o��e=���qפkx�t������]�o�O��V��f(�\z/�x�@P�p8��R��fU�j�nL�`v\�\fM����qY�cGr�?�������@�W����:��7[�zȏ����{�N�ND�v�bKT�
{���=��s,�{B-#+�Vx�Z�%��/�(?��9&s4]���5���3\>�P(y
�6*���+����&�sN}wT�$�8���/Aa�ԥ5i[����x@�� �`��������4�nc��,��R���1��q��a��­��[C���	�~n���7a�F��G�S̻1[�#ݹ rŀ�}�uNʂj*�6I�VU˕��UP�����h�1G�2�Rs���Ծ�y[�J�梵3d������A���i(Β�����~\@?�,�8�(ݙ"�i��ݤ�܇^��g�ms*$��ESפ�#-
!���U	�����lQ�̵��K�1u)�ױ~Q ���16������	���8@qY�&C��.:!�6��;c0߷s� ��g��"HSK�P
��10ڂ�|���}��([��`�d>�*��I6�c)<���H[Y�ғ���,~ �lvЧ%	Y�m�[��>+�8U�t�@�e@��v�AB�a������m����p��_ \�**�>j۪��q�E'|���s��}��)��Һ���w,���n�b*� M���1?VPg�>V{���M�|j�:`�@�������x��Ox6���Q���s5��I�a��P��'��C��ݽ��(��/(���Y�<x�̶H|�d��kѺ>�Y�G`���*"�r��l��$-.���A@<��E��u�#�n�����,�=�bB�B��^ͧځ[�<C��^� ��|�C$S+��G���.Ԟ�*��� AP�	�oe���W�\t ��i����� �D=CZ7��<���?��1����m!�����;ZЮ��|�-����;����ٱ��rO"���_�yF�
�`��!�;��U��X���t��(�JW9�~�#&�M���j�n �I=�x)��s�Y��rvHYF|>zBf�؉P�":�m��'(����n�?0 �捻Dr��Ox@{٭�Qh�BU��_FQ��(p��
�zk6=U�E��+��2p����v�)��Y��4`�n}��Ƕ��.E�Tes��q�e� p3I�k	Y�պ��ľ̫�}�Q�@�i���u��<��mЭ�6�e@x~_�"^X��$Ԥ����txY��&��_�/薳�q�1:z�3#9�Sd��V������#�����m8./����V+}����� ��jm�*~Ԉ`*P�,��\aK ������=}�������1�c,��s��E��J��3�2doR0�e��&��}
�)@h��}�G,;�`�͉BJ�Q��ib�]M%�%ᖝ�$�3���0f����9��.����l�O�u+6��,w\μ���� j";+k�Q@��7�HDi;w��d�N�Ž�͊�BX���+z���I��Ӎ�R��2��q�:�r��Ť ꛕ�4�J�\Dt��>w&�����Q�)�,m�k�b��	�KM�PA9A����C�T}�v�٥M���dҊ-"�Ҧ�^���o"�.��Jf���Q�^#��B6��&���(t�f�4��g~yŪ�Y5����A�Epq�3���Ĕ'�Д��*�AT:Vb��|���-%�uw�e�I��UU<��2Pl�SF�׋���t���ޝCɶ]+�7���Ld=>e�_�T{�+�F^Tx'M����DE�o�-l���P�G>���Ѐ]
�?�8a\I��$��B�Aِ�"�n��P�j�����Oy��eDH��t�k#�AX_�&��O�-���T`g��JK�7J��"�Ÿ�(64U��]'�YP��D���я���rZ~�xy���uu$|�2���d~���a�sa�w/���������&���5#k��'+��}PkH,h�d��v���Tϴz��Z��G�_ZN�ad$	c���Tx�4�nʤ��6�P�����ʞ���|�uxP�[�+l��VF�߃)��k�~1s��Q��"���c&�,�Ƶ�ͦ�X���ϠoC��l�I�v�$Fc�I��2!cY����RI����-䋴X�Za+K�k��Z��\�=�Y����n4a��gT���SQM����܁G�"�]������ ��wl�q-��/\y�u��f�ň7'�
�l6:�9��#�!X�Ě��b�����F����w�:N[h�[�n���=��C1;����M9"〧����;/Quu������� ��N�ۖ^$b����|7���V�Â��a��s�.X[�H��M�K/�evTv>�U۟��gSǄ�E�|���Hr2���}U{9��y,{�hh����y� h9��&5�Pg��X�s2� �b��ͼ�tzer��;�4O�+NfpE/�ݔ��(BW��r���9����(�oB6������픴Lq�K���xRtJ�?K((2�~^>��npM��Y��#�)a��ݡ"�#�|�a�*�*�j���[e�G(>�D/��(�|y�W^ x�m#�]���h��0T[fLL�j�~Ԅ�jo�u��9���p���r~��So��}�'�ť5^LP�1��
IJ�p�C2�����IJWC&� ���/��\���=%ݰ�){�����{8�ގIR�v
�Hp*Mi֪�X;����SAe���x$��V+<�$���s��\~�z�}x_a{�x{���#2'ͳRl"�/=?�z`��V��s����8�>�ȷ��k��*98��е��zy�i��S�h�4�?_�\;���Yմ%�V%��b?�����ܕɪq�ꑝLO�t���RT�^d.��p�*�> '����'b�CU/$mް�Q�ql�[�3@��pu��ToV�@���Wz$�jIgg.��]bT��$%
�?�H��4(eh��Խd�,�m��cn��B��
�b�9�uLT3��	yX��a�*O��;۬&����Ⱥ�6Kо�S��`�\�˙o�
��Z�d���%�����隲��/�@,���z��҈��I��cW��f�HЈc���h�|���Z#��Rt�Kj��N�\%�����n{(�ډ<��3�r��AI��֞��C����Gz�.Zm���J\i/��I��)�k|�c����l3	]݄K����'�q#��+��?_v}c�1N(��ߡ��~5�(5�T�Ӥ�O�!��n���0{HMWǥ<�����e��ؘ298���i���|IT�VDb�*y�>w����$�Om�~W�z�n�W(���r�
�z��Kȯ���'�q?Z�X���U/7���3c�n���e�����հ���e��Ym����� DQ� &5��}z)t�ȩԻK����k<�q<�2�1���<79��������8��в��u�F�'Z{r��(ഏ�,5O�o�ܙ�v�ʨ���Sn)ړ	h:ͽRj����D��j<s���Y�H�5R��z=�B���㼌��a�}���UZ�6�@d5�b��	��sV��5�n��7n�:�m��!�'u�	l��1*�Pte�
(���l��U��<$u�{�<l��F@�O���Wyl�@�+,�)����a�
e��k���O�X3��J{n6�Z���G�6o\�]ʚ>��R�,�g.����{Y��ma
/0���U�υWcnI�*%\��W�+�V�`õ�x�����b"�r�=�\����Kmk�)3��g3���	Y{�D�}<�76+7Ŭ柕� o�|feQFW�C�:?��\lS������[7tُ`@?����چ���� }zY��E=	)?YQQ��-ח�q��syBk�S�3Q�0�w����`�ӷ��FI�e�c�B�g�Y���_���x��l� ������l�MҦd� v��q�P�>@_�����^ZiE>�)>���K=��*�ڍI�t/��.%S�B@�����T ��/��GJ�{�fm^ͥy8��ro�Vö�ϿNo����i���ѓ׹F4�6�>jY�::�zֈ�K8�Ϩ]U5�SX��k�<����)�Q_���ߙ�%���sY���}�Q��*��4f�d�Q��*VE�z�5�
xI##:@�t�}��+�{�;��$Mr�J�������/�\��1x��U1y(¦}]ĤwD~���C���ڣ�1��H{�g�d��4=�Qa���M��QZ���ը��fGR�}�\��8Ғ�q��}�4;l��/LoF#�T��7����֍1�ޣ���'-�xT�C��h*��-'�I��M�ڈ�s��/�_�{�����G��L��z�����,�+����F*�޳V�����>S���D�Rg����;�m�.V<�����3�t�`#����N������M1��nܩ�7��u&�]�{جʦXO�k�௛:Rg�L2�4�Z��O�TS���q֟[� ���]�h���uj����X|��Vmwa�O��D�����K6}���n�Z��Oe��b�u��2��A�:vq��L�J�� C"<��Z��������������;��X���H���[���jB?�ݧ�#��Lr
���-T:�+�D֗��@�E�ѣģ�|Qgp=��F�uK�ܫN���Q��� B���Ƽe{\[7ҵ��H���n5֎6�~�b�.bצ�!�P�	�	G���k�눸������J�|������^B�^�Y�n����5��f]$g�(M,���D�h�t`&ȍ�f�j�7���xYg]�22X_7�����=��f��7*qKn�ֱhUr�Y�}$U��G�e��_~�T�1�;��j&�>��!��I�.�*۬�=��(��0T�	�GU�Weh�7bTQ=5�8�n��މh�\�_����+D��YZ�wr��V1Mw^im�G��@S�ɚ��� �w\E���Y�wStH���n�
H����v�.�ѥ�n�]Ux��D^����ї��ox�%��!�����NKx�#��:LۧYf<�0�W�z�4	ռ\agM�*�L��2�^caJˊ�:������Z�&���DS�zu`;%4��P���f�e�`�c�wH}�*6@v;���9_�ġ%�]���gƷF���S�T��0��o����� =^=�
���"�����P8� �ױ+^���#�3*d��T`� A���F�>�o�{�҅W=���ʾ�3�yq�z\�S�Ѩt����):/���G�*����fZ�5q^�3���XRg��X?��p�O����7p*�̄\���-��d[�P	M(�vQ���nS8�Z���j� 4!�f���&N!���[>��^������c���
��Er����ֻ����۠����q�c�]G�1}WUv仓!TE��d�*u��㴧����ag�1�Qz���,���R��yI�u�(֫�^�6_kk���	h<�"��Dk�y���'�ߋ�n�)�k�K�ngX,�h�{�]5Q{�q%��:�Dв��^ndH�P�m�R��
�>lB�D"�tf�����^O3�e�z�stX�g%����u�	��<�W<��m�Y� CDhkX�� ���fß�| An�G
�H��`�h"���L,���;/sC����HL��/�2mnM�� ��G2y�d�of��;���>$�����m=SfM;��&��n;	�,ů�)�Nl�]��3잡�.[;;˦��Ť��Φ=w�^��i^���`�#I������X$���}���L���l��4
��~Ti0�l8 z�Qٚ�(�~�y��H�`i2�>a�S��U.+׸��L��TO��<��u�@����#	�m�s��ӆ�u��*���~��fj�6���>�H+��m�8�B�������l==F���t��'Y����eo���|��$��tT
n���W�k#e��ND�\nB��.�l�,���=K?����p�|[��5��O �x5�L��z�L��Z˹H������ׁ�3�F�Q�Mr���4�4���2k���m)��4e0�$KufN���'W������L��3��̡���i��t��nQ�eJ-�X*\p.22�	`^c�9ν�z,p���ş Ɉn�}# 9|z!D�!J��W+�g(̏���\w��>�����	�O1���.��p���׹��\�h�(6�3��d'�jMk�XC�ݺKc�E���$K8s�1����m0�# �
�Cln�#z��gI@�gAЅ�t���:�g0��Z�2���	�1�6/L��%���I�(.-�}�g�
�)ޔ��}��_���OrV�^���xK(��Fe���^��"6�w9=��1�k�k/s�bQ�1L1ԃ<�)�N������uac?�{kQ���>��
@������R��m+q��j0ߕԓ���	&�Л�軣����b[`�����\�:��s	��G
�� q��H����r4K�;@��]	�D�Ӹ��$�����?�	W.@���)������%Eg��G&�Z�ɫv!%�h~�=p���~xjX��(�߲^0k����W��/	��kмj��P�
ʑ��Sv	�E��1~��R�)+L�
Y�� �P��E������=���WH�zq��{�3:k#� 
<.���?O��H�v���܍�M"r�I�c(��A�5�Ŕ����،�z٣�B5��~��tI��t��X�}�|N7pf���M�ڷ<fțP^�̙\}&�"׏L�p5
x�R�1yQBxV���v�T�%+�������j�n�	��E����#�}�z�-��S��G�=qN���P��76��2y�ɚ�����pQ�XW���4 ȤhS2P��+ZK��s؝ڛ��o�'���g����l~�`�f8)���>��z�����V��������?O��4��o��A�ΐ��&�d������^$�0��ٍ�47.V����9��B��OKH��<*S�����Gy�VJ��Eu8������\����)���kYp�<�l������'��|ݻ�NA~�ֿidC�量s�Tiy�E��r��x�?>W�F����N6a^����}̶Kn��
��-�����>��ݑ�O���ܡ~��3� �(��p85C���pR�n�{D*�Y�`e���zb�1�L���a�Z&�AE|�/Q�%н��]�d'�� �Vx���X����9ݵ/��t���n}"���%c�^�����u#}tD����@OK�IT���͛S�&��#7E�bή��>����գ�$?�o.��Y����DYP1Ёt��#��d �	�F�7�o�vؙ�s�5DZ��[ �w/�E�j�A�y����xR˚���cGe�����rO�I��d���r`�#��7�<Ʀ*Rv-:vE�ُ���?[��N�l�`0��_�����/�����4`0�Rp��3T�z*[�'�L�:��{e�]���z�	��*���I����ފ�j7b��~�_	���8�)��PV�z����D��8����Wdg1|�z� �(�߂]uB�p�:�%��dS8���Q�B?WE9Tt��̀	�ǋ�v��7��,Ö���ip@���ڷ��U�s�}sk���c���;���r�>l ʾ�����K2����"\ف�{>�!3 E���o�.����7��D��vv;��Zu�b�&(��_��eD�>2�H�TA�E#��s�"FhAb@j��%Bm�@�Yz��X��'hN2>��������M]����>�T����.��ʂ�`���<!`B�ju��`5r���`"��$	˔����T�F@�m�\�(k|����;c�XS�D*�}{�!ODC!�x1W`G����a�DG�z��B0�;�]�!� �q�F����?�8K�I��0͠����0�C�0\{�>�'@\�Cȕ��P?z]�*�1���e��C>@2e_���(U$���#S<0N,�t��i�;������'z��'�]�cDm
D��#+R���_Պ�����a^�����J9�
S��%t�p�������9�{�F�N�ǂ��;=�?����_E����g�Z=��;��4�2 ��)��\~����"36�(��C� G�)��T�pN�s��*?O�͂�rd�Л�_&Ϣ�{���vX�v@�;Iϻ�^��tP�����p�?�CG������+�D���o�s~����~ߩ�Y0�4��  Kn	�T ~} T��a��u��J��}Wn���NRVՓ�v��#]��9ʂd]�,Z���̭L Ț ������E��,�/�DM�/}j��HI�O1��س��m����N+?v˶	o�LQ��6�W��@\e�p��uZ2+7�&�����~!OV3�\�Q�c�0۴9����wN]C=��%2�N�b�|��ׂx;����t�E��4L�+��j�d6�YO+n�YUMP���ɜdD�=`` TΙ$(I D�5��^8њR���d�e�ɰ�}v߸п`Q��?��{t�LF�/��k5�Y�#b������&� �iw
:S���\�Q�vQ�a�(��Ͻ.�%�X�z\]��J�K4��}��<�ư*9��isx����?{�㕙* �(��z�׸��Us��:^��]V3�M�߼?�g�皖���rS���jjS�s�g$�e_2'o�G$�����I�w^��'Ӻoh�"��^��W0��rK##��9;y����܅,I� E�ӴMa�sv�!��?�t��� jG�7ښvD��΅�����t����s¼�0�������f�t�7��(}8�"�>�����7��fTP�Y���ٲ����A�T�t�]۪�pq�఑$JF@�@m�M����]��P�7��}���˽S��@O�!�ҵ��n�׹̈́K��X&)G�m?a�S�U#ah%��	��(��+������Gyw4�L7�E�;�r�\1W�}������Rԉ؋����R͚C}Ύ<���:<�����q�\����	�d
+I�~y�<xxQc�F�&	1j�6J¾�8���,r�z�]�U\Уv��.<�M�]���6�����I��B0�a,�[-�����C�o�0�qcè�����t���m��y��`r����l;[��j�7����_�:�����°ԝh��l�k�^;�� c�eIv��9�~}x=a�{R!w&��ݒ��b��v��gO�����\��:ټ�?�[Zڱ�i�	$H����;�\3G�s�k��"h��]3�oz�&@�NV�	B(����s8�WuM���؀zw��(eJ?����,͎ø�o�����1/�ʙNك���A�]>?��bby�H�������OYjŝ�.~M($k*���AD����9.Mn�w��sۭ;��WJ�u3�j�o���� �8]�Z��Ͳ�`�:��� �1H~kȃ���h�g~ã �m{�xJ�}���f�;_^ܽ��<k��>m�&p�h�������1SEi.Jƚ� |N��0� �#�i���_e����{+/"4jS��O;>��g����rAlP������/>àÛ�Rʓ�`��r=����*�U���G4��_fx�"�Ǳ\�X�A�9۱n�5���1��kЎ��y�-��9�1t��&�=�����hN;�}�.~7o�qU�+��照E&�V8W;Ͻ>{PB��ދ�z&'�������	���t���LgO
�,�9?{����@��`�7��������!���[�ʔ��H-20f#!)�99R�4]���IQ�T��f?� �o�3��>�%X0{�}�R�2�GK�W�5�l`o�AK�4H/����dwh�>-�)��o�C��.�r�C�f�����^�b��,9Gc{,^�9���9�u3����o���&�����j������-�T����،�=���t��������`�T����=q�����bff^���@�ԧ�m������_�ܱĂ���H���vr������=�q	7�Rg����_I�/-����|؛�>uɯ��BQ�o����Eþ�e�����A�!�;<�uz*}�wa�N�����&wr��?ȟи^�v��`��ԺP��͂�OB.�,r���	�߲���q��9�?;�Hs1��s��#�U�Ӌ��*��2�o
�n綱� �7g��J�-��u@M�q����"��ׄ�v����Ղ���vW�T�$������S���N�:~k�m��Tr��X?M��nU����a(��̅��o��i@��[����pj�rNpX��W��?�h�2�2-���`�W��/��*����؜Ps
�8 �� @��ݙ_�c���5�FL����;qA>� �k<~�Y屼�G���ōv�Y�7\/䃧�F�J�8O��.�Ҭ�w�;^���ӥ���64_�����
�Ƨ�g�l�N�]9�z�N$Pn�v6 ��ƤK�@���PZ�N����fM�*!��}]��`v����

 �)!���2CJ�����L���Ӭ�>��뭠7���;����@��egXa�3��ay4�w��)��/|)u�4��3��]`c4��<Iٰ|ԩ��T��Z�#�l���q���^�������<r�3{���;"��
Mw�����k���L�j{���i1ڕC�ch�3J6[�#Y�
�o�i�f�u�Z-�@���|�.�g2��L>�	����ʰX������HreA_�pw��[&�����_�{�Wq��pL{��U�w"��RMk����2�zœN<��>�4,M�z�B���~"�_�z|
j�l�T��Q����?{4�����~N�_�ƢE�v��H���ϩ�#��GO��M�/�֑�k�.H�s�>\s5��I�&ڇX�̒��g�0���u]^;��d:�����S�K@�#L�{�od�F�,H���c�\1sZ)5���u}�{B����L�5�?�T#^�:G�-z�u=�ь�FG�C����s�u��j샱�'��|��{���C���|���<$11��];����#Ъ��]4;�V}s|�f#���|НS��� ��m�J(���t55��E��8���K�=�)N&�}���U(�ׯ���w��(����;�%�RWu��J�Ś�I��~��KA��;OV�@�~>���TI9�cz ��*@���򈌴(��	������{��Ps%�n�E��轶g�;*$P��U9��5���_����wU������޲��*�w߬�P�D"��f��"��\v���i��T�ſ�D����'л�?�?�c����������!��*�r��Z۶�+����8�W��N4K����0��P�=A�Id$u�ߪ�-�S�y���m[�aT�����Kw��x_�ȷ��j�������hg����=���������7�0�4�1����@48�Iix��<$���1I��gb`/�V��R�l%��'�H%F���m��=����[��=N�\|��(��	/K���J��γkpۆ��ew���&��r�1�Z2���@`������lbj��/v>��y\m�@�J�0�,!�r*o��)<���QqaaÝ@	r_˦K�d���$�����k��m�=7�8�a��.ľ��S/�F+d�d��]���_���9K�9�ڼ�KO��D��sh�����=}|e[�K9{U��햲>���v���8�O�ʥl�U[�Hx���$��Y�/\��Y�$N����F�	}}P�!���==2�:h~]����y��cQU�ք+�5����LE礮ŭ���
�&3���O�R��u���`HUE����;��:(2S0���1�|�Z�RTW�[8{0M*���+Aj?���!nm�4��&��9���CO�ZF�v���|��.�^�kz=����V�ϰi��=�։R7�|�!hR�� �Ra,�7��&՞Q˺��.��#�vg}����2��B"4C��/�̵4�}�QֻXل��%oj�@�������h'$ЪX:p�¸�wh��	���t�'/e.83}���<.�;���8�U�z�������"���==���ӳ�?Β�:+���=u���oS/������U-���?ǳ{�)9����:}VL5�)���^��.��Y2ri�g1~��em/�{�ȅ }ȉ\�����ޤ����� ]g[�M��޹ժ��q��$�)]����(������)���0��j֧�Q~֟Y����A�yוGEwThe1/�67z�ظ�H�J(�''H��t~Ş*���Ҹ�ϰL�̐���!U��"�Y��f���g -����2���j̞�(�p��0��]���v�z؏X\���̫�=.�jk?��[W�V��o��C})M2_x٘��-����|1�<��JU��''�y����h�P�W�#��������bvM��e�����ְ��2~��N� ��M��F��ͩt����ʼ���F���U��y�\Xp	�Q��uչ�0Z�*�nԔ��;�!�k_��CN��x�E����PM���<��i�AՓ�"
����E����������^��7-�e��ƙd9ʇ*��x��JcJs�>�ԕ��M=�EC?x�#\I�g��3U�{7&��f=�Vwh� �l\l�h��t��+��
8��l�e��h&���7�<���)�'�Kf	����ːDz�r-m�C*d�dl�ou���"(�bV��_���d�#��a�4�`��O��%�lӑ�:
)����X�B*���������RN��
��sƁ��� x�)�+�����.G;�G���q�_����F�(���G�~��>�~_&�6��0`��(�[�\�N݂]\����t�?����s7^���//��s2�PK3��� ����C�FC���K+]�)��GCi�H��tG
���&O�ݕ�bֽ�:^��6�R����$�Ԇ�Ig�g���Q�ˣ�j�W�OX��W<�����DX|�����Uu���qu�	k�Je�Xpӕ9��)�d8
�Q�a�9"=g&���A4��wL�|���g!W�<�fJ����oh@|��|��N�`w�;{�>�r-W��nN�	�M"�}i67���#Uvß���+����eI�~�]�3}�eC �ؤ�qc5�
Z�:�z@��5(.�Ƥ}k�Zs����J�?1�7k����<�����xf�	����^���$U��.�Ս�7���7��q�gV�g����t��Mgߛz���j����Q�?:��������;l���0�l)�J@�@X��'��jwx��پ1`��p����~|�<�	>R-��鞬G�M$�_x�i휱g�i�
�7$ cE��ɸ~�O�T�L�I���o_����´�nI�y�/$J�L��ȆA����2�׿�F�GF�=�I	��a�_r˟ ��P��j��3��q�iL�N�����$��/r�J�o|���~��bMuuC��E���%�[�*R�{�����ĭ����c���όI����K ����u:�45��i㫴x���CM����8V/�,1 F(sa����j}W�I�{ZH@ڃ�NL��zxA'9��p���PJ���`|ĩ�֒�h���CO����t
ujL��Y�7�a����6�����w�o�x�3R��J;���t��h E׸���z���7�KX'�x��ڢ�ULW������ipw���x�M����^]��;:E1�b3�6��t�'�OB[�0B_�i�6���,���Y.L��y�ܙ�F�ouZw��O,3$m�r�}��6�>Cx#��t��8�����QM/_ߨ�c��X�
�DzWi
�;��^#��HWz�{�� ��.%AZ(!�����9�G|����u׻�k=�יٳg�ޟ�e&|gB�/�!�>��	[�^l�I��۔��<$� ��rŒǅx
-V�-��T����T��h9�	��oXi�&��I"���yEH�;~�.k��b��MԊ.l��d���u]���m
��3�����8'	�Z�s^eh�����<9�hW�!j�S�w+GǪm����o���%��#*��x�������i�]Sr�ytfh<Y]�4��i?O�R�/h�7�$]��ث�f��\W�=?.-3Z�X��e�.5���'��8�o���7�zj�3_��g�E-S�a:k;�o�3]�Q�j�����������&�y�b�kJ�:%�h�R>��9�!j�+���� r�)��(�8}�S�۸np	�}-�hI� RT�L� ���<���fH��n����``դ�+�r��E1l<��
B���LrB����G��X�c�[Hd��<6�� �/o�M�R7.u�����qt�i��ǰs�3��\��h�#��ʇ�]�k��|~;�L��y`�0'�D#�L��J�""*��#r��6)�^!k
�����`O�Y�0�m�[����Z	>'�g���])7)I��\��6��*��8jO�SjB�6�ȨUW�m���Z�=��6-g��X4OK��K!i��@mx��=��:@����"r��CE��"��i23n��FƬH�S�U�Ca���m���Nc9R�i��,2�Rk�4>�y&���H��^�OR��cl;���*Z
��Y���\��&7�X�s�@��w���Yw�~ W�Wǵ:���E�B2�s������m��#��jz�}���rV)�|+I�յ�y� ���7&06�5}O�U��/�a�+�~�b�m_ �f'(��޵_i�OR\n�@`K��p����>�ACf�d�<�j�wgC�_���B�)��6�ͯ�ne N��_�FA�sRG�{ô��� >Qį����U��:s�zOp����551y����8́�����G�������.�k�5o&���(�Ɖ&dd���F+�q�=�Y�"L_�G"2,�T�嚡�'��ܵ���)p�`��p*o�C�EB|s>>���!}t�挿����qZ �\���mK�W�G)��|s�Ɨ����s��k��s_���d��#�B7�1�
lBR�EH�u
�|���ǝ�Qe���%�Ñ�u���J��%͸�4��O������~�"�͢����#0�OHK�ǃā�8�ǀ^�B!}S��F����Ȭ݈��j�ykG{�A�P㞣x
�o�USu�Q�[��ټ��!�
e�T7f�<bM�īvk��ZȦ׀�Ɇ�j�$2��N��&��ϛTCۻ��o�&�k/���u6���[,���6!�2BjK���x@�轅+�,;�2ʻ�n���úL��ب���:O�Yq���5��+]}�0�b>M�[��V5*VRɄ/���ARՈ��o	��<�v:|���`ϰ^Z�ƹ�I�C���ܝ�:�TY�$t�Qr)��}�jM��CTS�k���v�1�諸�[�b��nv�;VQ�resK]�\n�dG����'p�b�V�L����k��m��_���[n]4Wh�gGi8�"RW�h�n�ʷ�!���Ş�$�3�n�w�-��"'��4��o�	�YWB�H��#�3h�D��_�mA.���9̳%��q�Cb���{����Xrz<B��f!��E��[+tX�z�(P�rZ�`��z��*68���E�m�NY&����n��<a}�(�j��Od]KA�vN�>�e���+]�
s���'*vP+�>	�-�6
�[d[��Yj��oh�*�кT�:z;�38߲� ���ƒ�8k�vW�7g��[�7B%�c-���M�M,�*�q�L��.$��$�w�?���=a�Q���5)�$�
ۋҰڞ�}��s���lU���^Dg)Ќt�q���[��������)�&�>��K���6��FrY�`{|QU����=�20
 �*6>��$�O0=�U�Mbّ��L1%ios�<p��l���ot6�m���oI��V3b�xҠ���W��Ob����A未c�[��zq��8$�����:Ӭ��\�o��Bܠ�z'|���I��zẶ��[��5D�k��+��
�J�'W4�����yߚjYE�l�%6΂��{#��+�_#�{�?�9���X ��}�U���n>g��͕�x��C���Z�~�9��ۮ������DX;h7��wH���~�@@��d:t���@��%�P���i�Z�HLLY<su����u	�⮦1���}qa<o�x�9�e�?n_�|�RQ�
�gT�>�g9z����j)@m�T�V�]�l/&�~�r.�*�A�{#w�dլ|�:D��+��T\}!��³���#j��� `��:�$k�ڎ��>0$�<@s�[�9}q
�K5M��$�y���"�'�k�Z���E��M��|c��:��+w�e�@�a|�;l���V擖�:]X�b>TVw/�2{��)��5ta��U����.�k�3��w<���ٓ�ҜD�1$��σVk���k����-�{������#h��6�ŝ��LqVuSU�`kN{�嚰_�M�.��}�@}��ul���Li�S��g���5]�+�-��`YTu��x2.��e�̐hY2�~�=�j(���UU-�7�&|����Z�"[�%���dt��W%Me$��ɒg>|��U}Q���h��{�=�4G_��x%�1�w�^��R�Wy�[�̩h�h��B�[�B�U�r���Dҝ͞��V��-0"(vߍ��X|�����*���*�l�DS���d��Ed�L�[�~G;�f�Z-�ж�%�Ȁ�|�>�~�@��Lh彈��6z��Ͻ&	e��J� LOot�:x��Zg�Ϟ#��(#���.�Y�L[� kC�ի�.������|�륟���a5m^�:V��Q�T�c. ���X�	�BϹȂ�fe����99
/���YZ�h�c���Щ��A�ac�fӢ���ojA�_�b͏��������ߞ_ ��z��I���:/ r}�,��C "l!w,d�{q|��Ǟ�������sVα�m>�Z�D[�N�85�
�m<Q����)w�������C^EnQ�S�w2��X�D+��J��0�Ub� ���Ė�S��r!-f�X:m|×/��R9���7ƽ�4u���]�&�/i���Ѵ�>�`�rX��,�,����q�ߏ�����jk�4�������$S�t�Œ�����o@$�q-��L�`6�L��Aig���gc�ᶂ��p9f���:�����F�i��}|�.��E��+�ɴ��[}�!�377!V�W��v� ����(���fūj1��i!S��w�x�=x<)���!5����~U���)Db�[f�:S�i�4�+Ͱep[5MS-[f;�/-�4�S�mX�g���e�8��E�nIV�߶��<�IR�D�+��s�
H��ZU0���Q�㙹��%*�D�r����-���G���w�����׊h����a��-R�U ^z/�_-�]y�e�8;�M���+_S7B�4�
���Ro�y�m�+?	����\�ݫD*�_��&���NI)�;t��&yñ][+�"թ�!y��˙�z�Ֆ$YC���0�e��[|ح1ʽ�y��OM�zܭ��|q����VΦ{U�Ѻ�z��֘��XS��y�"|��;�i�x c&3�ڷ��k �Oi��[ׯ�6�m3=?�U4�ݴu��x��#1�x()=ׅ7��'��B� ���Y��idr`�X�oH����5�2��=K�hla�h�l��MY�^��$�N������Y����*�� �R+����-;��ؕ����kƱ��[9���{o�XV(����P0O~����NV c����r��S�E��"�6���@����w��Z݁�#"]�b���)�(RazG-�UC��gp]�9%�dw�r^)6tt��pҷ� �7��uX��g)k�5��q�x��G�
���6����^K���x��0�c�sQ�&�H����a'�7{R;���l?��X/����
Q�^*ik�����8a^s<e�" ��N��-�9�t��u��!P-�����'�CAէ�W&�r�+��f��]�߇%&a�k>���>֯�����JW���U��Io�� ��^�������޺�ni�o��t�_T�u7-����C�$�H�l�7w`�k����Q0 S�[�f��~��I�\��Q��'�6���L[͕6eE���*�#��	Q���3�R?ې�Q��"4[�3����ʘ�Z���eM"��\����.�4�\E��s;Q�i~�%X��X��@�G��?�9e#�~ �N�DV����X��&;a���L�)��6� b���w�9�����:��>z��w��7���C�5�&_@�	iI۪�|���F=��lG�2R޾�wyJˑ�{{�̱O�_U�S$z�3�O�qЫ���{���E*#1�x���P$G����GƄ� 5�M�'�<��|����9�SLf)�Dn.@K�׬�D7o�Љ_��6`6�^w Չ�� �2�+� �D4��(�^�m������@�᯼E�'��C�șq��d�Ze����D��]�.�+����:�t��ʐ�5�>�M�w;+'v�pX�<9O�������r-nst�o�Ho�P�����ֿ�<�H�LW��Z�eN2��4���O����ؕ?�{?�id���;�9t5|�0��M����'!�O~���ᰣ�	����E�>����)c
KV�z=��v�cv4Qm�]�%l{_�/���J�z�DԲ%�������T:�G�� ǂ��-�k�=p
�h*_.cr)���b���n��B�����M����ŝ�@7wT�
�*�u}��ļ�>�Hnd�m-��t�S˔`��mX���?'[ǭA�64�3Q�E��u8Έ~t5xխk-h�3��	���f>�9�r��i���t�m�W��x(��;N��&���C�ig�L�K�yeMHJ�7+<��T�I�������U���o�,���[U���@l{�zh_+��~��y\T{�Z|
AA��S$:w��	!�YUa�|�u��C�^U�Ms�����Z�Pqc9c��V�/�a)�
�~�F<|'�6%�jk�)��@��v��x����6�E��EK��+�rx��u|PH�	Qq򉶵�{�T����O�ԽOڵ\pL�Ś�%��S}��pKqE����'	U��8VP�s0��\:�T��5�(<��'�K�Ι���5.�������"��U\��H��"N>X2��f�p
[�e9� OF��4�(ܴ��ͼ���)��t2a���(��R]��*�
�2y B�0�,�
�I/�{_/��bsw�y���??~�U[a%�3`+��կ�DU��ǧ����>��1Q\��
�l�����<#u桅'�G��3�������@��:�[��Q���a��N��м}�Ĺ�*���&W,���.�8Җ|�t����%U�Bk;ij��gpM�̅�v!)�\o�g*���bm#I����a������P�!;�X��Qvn3OU�L<;���tENe�[�@fv�p �%��s=yd��ѥ�~��]�]ҹ��N��k<YZ��Tl��c1���1e���\@YL�Pop�R �[� *�솆C�XS"��R�O'� +?/��$���U����N�z詡����-�Ƀ�-������y�z ��`o w�ne����~s�>���2��Д����R��+K�M��]��tų�Ӽ�%(ķ,a���5)n>5ޣˡM���	>��4���;��N���R���2��R��&�b`�\� r,s�����e�$��D2�ɑ���jUG���{i���XOmu��[���T܋�3V��%_ҝJ^�:K�2�����ƻٳ�P;\�~ϔG�)�Н �|���R�����m��r��[W꼟�Fi���ɯ�6�|�^�^ee�Ʈ�trL~'�݀���ee؉)e%�X�����u{}N��:�!��l�4��n�c���b�܉m�?��CN֖̂Qq�?��@�^>�f�&�ȃ�[o��M�B��M�"xj�O���l�=�������ǣո��x
�iǩ8��|��s���׶8iw��L|_u\�����c�"��il�1�>?�*5O6O�@�����H%r��M|P�6n;o���-8�BK%_	I=~܋�ۂ@HSVAeU�LV�򛊷�y��t���=ҫ� ;_p^y�T)|Y-ϻ����\4!>��z�B.�|��҅�<3{z��Psv��Y[�Ϗ� �L�6b'b��:ې�싮�,����=���7�$��,'�1w$ׅ����C��6
@�9�J���F%Bt]u�*�+���4�#@��߿t��*0�iZ��!a��I�VjOc�т�qq�K|9��'�Q.4Wڐp�~���D��9�I�)�y��N�
Iic��  �A!��n I�p�`�p��[q��9���6�HV��`�WF|	AVMw��/��H� �QTJ@�˶+�Zt��5�f׾�y����8	;`��H|���a�zk����'ʧ처�S�v �Z?fIﭠ�1��k� �X!��e����^c(D����ߊ�y�E�A������F���)%*J�H~DR����K�I�,ѢU��A��;a���j�]��-� �0��6�%���YEb=xk��5�Bt�h�$��R C9���N�����ҧ���&Egc�)��7�:�(uaU/(=�H)<�ꂊl�\^����L�D��JS�G*!��Թ����6�U��O63T�����R�W��NIt�z�sڱk�`0�-3	 N�1y�S����3�"�꽡Bg�B><4�d{�$	+b�Xez���zԞ$@�	K��2���9�:\d^_�݃"�u,Օ��n�UV��Rd9��s`6w9[�� g�?l���R��c� �h���cB�b�������^��*�q��9N���*vLZ�������e"	�أ��Kޱ��$Ia*g%��.��9���mXj���/�1�j��@p��d�f񑈂�dʗ�X�S:�l�.f�w�e�u2�߾�dr�}�<(��1���k�}��sJ�Xm�̩J�.��`�GGr�ԉ��@����]3��������^LG�e��O�2G�n�"�� �7��aʬ�ry��7�ۼ��}b!�����Ĕ��e7�WW�Uq{�H9)�ޤ����O�b�G�x�T-�gK�'Bh%j�2��>i�����ȴ�cJ�/De0[3���c���p��'����ȳ�N��&���%H�o���3s�u4)9}|�=�*�,qV����߲{�+�[���_�L��XGY����d�m�nz�ƽ��%U��2�Yʹ���c%$��Y"������C�=�`���Hy��*�C���@���s*R��CDÉ���Д4��� ��9|�)��׿'I�.���/�g�}1���������,����j������ ������~������I����w^b�����^����?#���S�Bw`�������86�L�C���0����^���%���|q���9=d�4�+�ލ�l��!��]�dϮ�Y��5�:���-����%@@f[�J��'����@`�Z4o�k8gԋO��>�F��$_Uy��D����L���o�soߤ)Qˍ�1k�T*���Qd~����'��<����c&%>�:�=*�k�-�2[V�z�>�f^���4}'Xh%�3���Ĺg�X��~�~0J��d���po޶�ŉF&)�CZ�&�'H��JP}�<��f�*'ihV�����w���D�2����}����C�AA���Z��U���{�3��߭2f_�N����7P#:\�`�[�Z�ïa�8�}�+� ڟ�*��Y?���pMv_)��2�Gz5Ri6��t���:v1^�^D��lk��Z��$Iվ�WJ�܌�v^K��%li����~\�x㓈�v���(�!�8���w;�E�&�T�������
����Z�+���^��s�c�z�A�Zk���[UM{�����{�a~U}	�g�0|���RH��^��� A�|$�x�*�Aά�����"vW�n}#��r$Q����@v�&�4�[{���Y�غL����M`���Q$�|xq�xR���#l��#J6nf���̪�J����7�V��g{"���@��}�-|*�&	��|�y��
8����s6�����e2%��
����X��C��}�U{�T��
khO��
1���C����9�p��
^����:ع4O(�mJ�A��g���!���{���+�M3��fP�w�&�OG?�|E{Y(B5\m�l[��'��l����Zo�ը��
�����aJâ��K�M&5�-,��H���md���<�j||>"�>_�T�r����~Iq����[�}��Hy�(TM&�`��i��rGn�t����,/2R��!c�V���{��{��۲N�ǈ�@6p��&���z�F߷ �=���!i������S�c�2!��C�%Ȃ��;z�b��c@6X�=�j�ve8����4i�2sF�೩����(��"C�À����a���`�����pn�NV�H�p��C�FDD�33Ծ���h��AO��+��e�&���ѓ�)��|ȉ�B�rOxC?��D�����9@��햎ײ6��c'��y(9�a�v�hV�黎�X4d�j�;�����+�v�T�����8�#Q��d<���õ���-��C��&���cD\D��O2�����+�`��J�VP@�́��Z��!��6�juu���>-GkX.&ᙑ��0�hw�¼TRp��W �W���u{
,>MaB$i�R;2rr�Za岦HUϖ� 6r���-Y�tH�;+�e!�������wH�@��P��|V#kV�ݬrO&1���8�ٺ�Iص��$���?���o�lg�I��D>d"���L����hM�b�(˚{
���ha�\Z4\{�*4�@n����k��i�o.���8	[�t<��q�(C�6"��T[$��$�d�~6<��RL�(��Ob��)��\ �J�]CB9��e���n��,��4Rqp�b����gٿ���T�=C���i��{�l	�Qv?��Ņ�W��r_�C5��;�K��V4���0�ј�[�﷏�=�[�٪�����ǻ�Ʋ�~=y�]�9-]ћ��f��f�i�̺!�	�b�E�����(w햾�w�Oy�_iٵjﾹ;)���}|��8jt�Qvɦ-� �����OD�����gt�m���'�䞻����!'ݭ��ok���W��Z�N��}k�L|k6' ϻ��~�����銿P?v<j�J����?k��vtH���J��x��*D���E��.r_+^�����D���+���$��[f�;SvW����J����t���5�����U.j�	' �nw"6�@�����0�W���,�+>
2��씎E������	���QI���0��>�ik�N,��U#���p��r�p�ũ�V�}����o�������� 'q����,����6�kLW'rx��e�>'Q�u��j�����S֛��������a �7��
�t�Y#>��#�5}Oj!غ����ݨ*�*%8�U@Yp�έ�njg�ԝW���a�q1QG{/�-0'D��������/�������L�/�V7=^�{:��R����v�cJ�h|���\G�,���SSo��*��Y���d}���iX����wT��&�0��M����� ��U���jq�6eA�����|�H���B����� ������!<.���@\�j-$��%�^�9�M᫴/T ���ơ��;�}Z�Eҋ�V�9Mm��և��ߤ������TdDT����i�0��9�(�U���YH\p�f�ïL�<��,�����NU�1�bg�>�!�7�W��8~[��!҅���<o����}O��А�]�������i'����:=2��m�^�=�E���4;��z=W����t}���B��#��%Mb+��k|ޡ���	��@�PuZ�l�ע+Wv�y\�eWf0���:u�i��b*p�}={|2$ry�2_�ʊ��7���5��1��&�ۯ�����uK;���|5�=y��4�5x�B��]T��y�(B~TOA8��6���$N�p�ˬj@ZyvHh��jrM(b���i�>����(���-kr�TŖ�����u��Ğ��*��z}��k�6� ]	K�~Ř��p������=�.O(��~�[��Z�����\Ӣ/́��/�ii��yը����O��%�[A?�H�>��䞿N�%�8&�IW��ү~m�Sǁ/���ܤz��qG�Y�,Y�n��ք�zD�!�����e>+P��vʫ�~�=������T_�e�>��|�wJ�"��z`�T�+�;Ojգk<ޱ&�]o�Ђ싮&Z�2Y����D���)j6��p,*��֏�|(�@���E�?��M_�[ �*\����缋��zE
N6���s)1��6J�6�������rDG,���x��Y�Jջ��iЂ��B�|n�E����2��4,�iN�Ep�݌ii���T1҅T`���]���W *����oUS����ʆ`��<X����3 Xx�b�@�!�7�\����!�!�4��3T��hF�Չ�bx��M�}���i�K��+��
���<i⦛I6NCwz��m�v�F#�R�r��5����y}ҥ���7��N`�*��½���s�O���3Z{7+-��8��ֆ�V��Y��7<�i^��;�4eP�a�hi2�2���ᕧ���~J���<O��%�Q����%M`�ƣ'��9c��)�.Þ��Z�*NÞӒ���g�6D��z殍�:;b3�ӊ������n�e�秫����\N�`�9��������<v7���Ƈ�$~o�y���ޢ�:�0g�y�%0�w�Ea��9�^伛��a,�M���;���P�T�)�3l�%���q�>�S�߽ݱ�������]��'�?�)�g26�7���`���D<+.��ۏ�?��L����)���DN3�����79��<�ʜ��%�pjʤuֵ����	=�n}����M�S>�O5'���k�1v�[Ke�vkS�.�����ݺ�)(,l�1�����h�5',q\�MgX!U@�Ĭ���5(��{m���W����9uSS�A��������k�r	X���A>�<+�U@��tБ��=���̵Y�WB[͛�$<K����EL?ui]̺Ӝr-f����w|��*��>W'V5?>%��c�F����LR�u��4ۍTa;Af���G���*��n:�R¹/�|���8������[`u��$�-���,�������ӞZ�0_���� �RH����sԲ<�<���GaR@��y��+	�Wn�?�ʜ����%h�!��(�l.O~��Z��=�*�DI�]:�S�G�`���Nd��������kVb�&gm� ����'Y=�hO{Ƽ��}���N�X���
�����[�\�����?t}�V�M�0C���o�\'�>�P�?��d�Qʨ����1�y�[�)G���j�n��8jf���z&�Q�ityr#�Ϯ;@��IׇV���\�|ˉ
�|!�$"BWɱ.׆(Y�Y;+/�x������^���z2�U9�V;��m͸ں���Z��+�Y��8��>��-T\^��T��Џ�䝒cq��R��m�\�/�5a[]��m,lEJ��Y�Э�4�9�ǲ���c(����_Y��[�d����B�}v{�x�f��?���Q�������r��FW����䙩��r��`8�礭��kK
=��t'x���-�p���Q'</�+))Io��N���O�b��A/]����j'l>�^s����Jٔ�hy�ONӽ�g����ya�f��A�C����'<�.�� �Eq茈���O�/ӎ���%i���63�����e�c�~}o�>ͩ__���i&F<���W��i�;��ӽ��J�u}�6��Ox�衉L�n}���>Gu��(g�ޝ��[�O�D73�jڇ�����?��L9l`N�~���@�J���Ldtt�#�^)��� ���`ϵ��G����՘A�{~�]i����z{��3ix�U<1ES#{Ү��Օz�E�i$G�׉j��5��ΏlG��� ���QZ���B�]�Q}�~��Դ]4bc��X�s�����JK)X�y�ݑ4ϬfEۈh���Z� k�iJ0��6+J�~��I9�3�1����)������E��(�ds!F���pv�쌘5���^���y˹��4V@��f�b��#\�~mmm�di.��$E��/��;i~dH�'���kЍ�&��K`0��Ȅ��$v`T9������iJ�w���]nz��?�9�iv}�c_D#�#��� �:�����N�>���L��c8���Xdd�ܑe>�<k���MrV������P�;�݇�9z��`�Vs�P*�ƳcQ��=;;޾�5�y�.�;9bؔs�ڵkĦ)^>>#E£iJ���-����BQ)�T��Shcy����]�X�&L8��M����P�@�k�#��������QUMmֳ�d컿�q�<1������5S_jSߍ�_���@��5���1��!�6+�MS^�!�V����f�L$f�/uf��)�n�a��]�_`5ݹ��3�4P���:&s��۞$�#�7;e��t�5��\���gmy5�5k��$Tf"�C�'ݺ/�w�^\�|j����K��5-�*R�@�7ä#n,J�����p�NJ��� (l �!�TU	w�^7�t�KH`��l�%9��_?;#�+ ?6��N��g�Nv����u4����e�d ����uj#t�jCG�l
]hQ�A��陘�\io>0�244�Ƹ�O����t��ׇ�\�Ħ53X���1���dB��8c�O3��,�ç M���K�����0B@�!��R�GA��۪|Ǧ�� ��T��$�۲�w�G&� @Q�m�!D��N�.�y�Λv:���`0M۵��ݑ������@+��6�e�7f�SRRz�R�(�Gp���L䔖���!��e���?��F������FH<�i�|�y��n�%�,/�.�y��1C�-kdj�/x�HR�ABH+q2�;��}]A�f��<�:_���jW�/s 	hӯ�B߾���<ӛ,�ׇ?و>�ݞ@�_E�n���^�1����E4탊t
�O9�`�m�h4xm0n��]q�{�`聑��z穆`��mf8X��w����!t�;ݦk�w5�1?7�K��������"�[�SJuL���#�c4f��C���0W@� u��y�ޞ��Q~%�X9�!�~��+°�gv�k8T��y��<�"�i��xe��z����i~��>)""bfq�������ג$���`������?��������Z�ciP�a�-jj��s����Hg�b�e�8��4�d�FW��ו��Wk
��.N֗���</�{7���B��<�#[��wt���r�4�Hp�~oy��Yb��)\s Ja����a�!��K'�!�F!��ԿkN5��5��f9�~���fW�A�B����;�q��4��#���5�%��y�ɺ���ݼۍ������,.l��m����Gwc.ǜ�>J|� ����̧O�0U=����NN �0ź��Ͱ�wu��n��������i�����\j�+�9?���ܻ��.o�P�>|k��33\�~��S#kQ#���ܝ����@��XǫS��aL�!��g�ai��U4B�	��e�c>l�1|I�N�X����7�1}!�ߩ��s�{�������xえ��ʭ@w��&��-H�w����[I���΁?����.��~���j~9�k�_�\/�:�Fs Q�#{l���3���.����us��=dJ���J��á��GVN�WjD����"��O�?ן
=�ރ�0�a(P
Ŭ�f4�72u��F��4�,s6oJ�(�j�� G\�%աV$5�cI�'�;�� �#��A��i1�[_Hc��G�N�`6�N�W�68���!�� [�q[��Ą[� U0���s�Y﮻3��̑�3^ 7X8�:|bpp0P��� `�����fA̛f��/.��{_G�����:��*ۀRpv������	O/��A"1t�]��JO�ز]��׵�k#�#]�ă��*�@f��� �6�0��U�u�FĕK���~7����y��0`��r�գ�-��uu�&N���l�T���B����>bȄ;����*�s7���s�K-�#�K}H���V3E�B�w�q2�1��o�\��^�4:qFu�R�̐V��iAd2���%�.|p���S��[�}����AT��Lp�]�#!��5*��pM��Xp����#�rt�$���Z5~��>�	w�e���C�B>�(y�i���|�ږ�C��ߵ?y��[�D�`�(5�"��i;ފ��̯�@j6��i��V
��_鵌�Z�o�d�{W�<~���E�#h�l��$�\jTS�8ɥ���Lpв/����s�QGBنPQ�EA��7!�����k�ZD�+B-�f�c`޸��t�"o�T����'T#8>�F�
����W8S�����([U�F 8J������k<�o'�n`�����3��kߍV4B�Y鎬��ݻ�o��A��7��N�T-�F6���g��PB.;�*��J9�+r�/��yF����X��8���zn�T���G<�QA�a���ܩ�a��^��,��
v��/��sFiՇH���s��>�q�'+l�J|�1�d������B�xvv�DyVPa�R�e�0���6m���M]<uȱ4J�c���X���ɽ�eUs�dnGAv����p�� �R����9E��z����fEw�W�@��.�1� !6I��b!�HH�R����5.h��K�0;���1�wO�"À0����N�s&�1��5�F]�Y��Ai,�Xƨ���2�ʉZd�&F;{^���}iuv�{s�3Fri�?r0rf��$H[�0ȌX�D+O�;�B{��#�6[3�x����V:�@�Vz� ��:��X0�r��2��'��
˄*{Њf�x��	O�gb�N���O�t���7^~f��B�|���l��o����D�*�R����l��/�gEWk$��r� t�OL��˭�9����i�w\jN�\ҫPS�4�*��6y�`��CM?ɛi,B%$� ��j���oȥf�@���x3���#�;�Ԝ0�A-�.A'#f�VWW�b+���m& pU)�rt���f�I5�yp�<@r����� P�O[m�un�D��v����$�Ù����v�����*�I���f- H��v�Gieq�(�xfZ�8��ˠE��w?�a��0�������/�������C������xV���X���R)oeH�D���>�7�D�ĿI �f�������B�P�_��kte����
(��M ˰���#<ѵO���Ȉ)
~ix��7�]�]��a=�p��������ֶ8�wx��r���QGy���/S��	eh���TR�_���,��@��@�u��31a��~Y}���'p�w�^�����`C3ޕ�~gL�swt�%5�H3gۦ"��2����܎G��.�|��?�.��`�/�A,I[�z�4��eʯ1�+�s����8WY�Ɵ���IE������	�i��+�R��p�6y���N�Ǌ97�Šo9����!<I4bsrA��+h]k:
��5K��J�L�S����:�y|�PF���O?�mɓ�X����_�'���yY�/�mG*� ���$�d�T�p��d4��?(�%�nx,��)�+)� �o�G��d�F�E����;��[�*#���s�L�~.�%���lu}eBr3�>�t�n�h�z�pt��Ȧb�vK8N�`�2<��F��3���eƺK�d�te����6?�س����{�G�7��e i��x�r��椄��Q��$(��P�}>IS���%�'����� 	A��Ί'R�q��3G�`϶5N�bHT"�	��PWJ��A�/�RM��G����EN������
ZX�X�^�i�_ڒ��`�s�\U� ��Dg����B���3�&��&�0�+c�v��\BQ�v�`|���Y3�_�4�ܴ:�s��]��/��iǀ���|^瀚���)p3�!����_�T����_��_2Pל��z�+��?A�_�����s���1j@��?~�e}!j�B�GG��$��?Ww�O���i����E:������6}�:�ԔRO�޺����ڰY$Q�8W͘)���J;s��٢��SCr��z�h*G��@��������V����{q�j�.,��ڤ��࠺G*�j���[�>��ͭ,�V��&#��C����)�;Cھ�OteJ[���D�C�#�#I�LD~����������w���Sh���ƛ���d]kh��
�׈���F�֫�5:?���&�4���&�E�ѕ���W�]1g�hҢ���}�-�(3�#�kلL��`H�U�ss$��yh6�j��[J�~ֵ	9V�[���f�O�'�O��K���eX��Z.��ҒJn�_ɤ��aF�8C��M��@��4� �n���7��}]�]����$4S;h����Eú��]�5��_JF+�90��r�:r�͚:���s�Ṕ�T���
�l�j��}v2�ݻK����\3 9"4�u�ɝ�\:E~s$Ƨ�}P�>��K]�������2�,�+̻�a�S�ow�rG$O[^q��_0�t�|��k��ނ���'1w�'�row��H:�f{M�U:W�ƅ�"'w�;H�֜���7vp�mR�S%bg�y���J�;�rJ�y�'��6&�]�:�{�ѧi��{D��azU�Z �yb�ۃ�:����'C�[�8~ћv�Unx�Nϣ۠c��_w��s�=/��r
7���gs.����PMfQ��#��)�FP�)�;
�(D��4�HE�A:""-(ꠔP(]�H'�z �$�������]�w_����Y�q��s�>���v���\lUu��n����p�e��^�i�kWJn�b��4-��/z:����{�y���hK���q&�j��|�{G����e@5���mR���ni�q"n?~pb+��cV
4��� ���58�w�����Tg�ON�-@nn�Ȕpt�hB2�>Ι��^�m�c:���f��n�x kr��6��M��{��n.���]��	�^��;����w4������(����?�D��O�?�D��O����Q,w�}��t��������G*�a�j��8��ess3������.S>�.�6��E �M5;ח�fw��<G}����
,�KD�r�䕏(V�M]wi:��Qz˽�w�ƈ[��N�}�<��HS��ȃ$�Ra����
@:e�I.����x���pj��E.����͔p�4(ES,w�5>5S���_��Q��թ.��:�q�d����*�]�O��_���(��.��k��B=�!���|U��5B(��t�X���n9,�U�P�0��f�O���Fn��g�WW%����{��}n����W¹��~��O�
K�����=>����V^<�${�n�۷o��~5�T�P��RI-��um���dP��k��9c�4qM�;y��^H�/^��@��gyp��2��Í�Ύ��ן����.���<��}a��dT�_�)/]�F�r��)D��oom�ඬBH��<QUES ��HҾ���k �=��q����;Z��j�[m�;F�����	e�=��%-�g��V@yG��*�_�П"���'��FH	���\�t�α�[�Ł�2���<K���w���~���'kO�	��Úl�p������Y{T��2tJ���H������\$!g�7v���1�����#�#45��^��@�!�j�5ߏ�Z��A��0z�֤�hȔ`��LW����`���!Ͽ�0O��No0�65���]L��X�ʽ�&?���ի��mi�j�,� ޣ���D�%ni�H�!��r�cD�`4)A�љ�<��n�����3�a7l��(pUY��u�8��"qi9��bBi;m���IF֖�J�?�)�:�G�G�r ��sjϏ.�˯΅���\��2A�i� �咱��&�=����DG���1��_�V�yɸh�;�<D�x��y����It�����0�#��xM,_D�*t)�f�K7op}�%�q���a����m:6|
��1
����
�?z��Z���!G��l�y��,��b+><q���@\}D /}��~4���1:\ӟ�}��h��?rZ)��u��4g�����u)Z_M�zN��; �E~>-qͪ0�>u^X�M�M���Z�l�%&�ż^[��lME�Ѫ��PNvRMJ#�F*[ :#'Kp�?��yq���l��g���$4�1�fu̪��*������N����T�ՠ�'�k���u2�د����[#����jl6��p��+���u�ܕ�A��Q��oȺ���E��L�����?o��JQ�BQ�ZG�
�[�UK�]S��#2���H�����x<�.�8�5d]��{���
�zN
�覻o�����\*0pjE�}�@v��}c R?W��w-�p��v��8pbǥ�};�����������_��y�����/�<k��!��`-���Y�l��dԗT�������{�\�דN׾���6Ɂ����YJ�vk?>HG��sg �0yQn��k�4F$�5Į�b�Gx��U u$H�>�]�k��`�<�c�b/o�D]�^�����7f���������1?(|�:�N2����1��wא��{'جn4��>R�:��#�<f���L*|ϒ5�x@V��Q�k/%4�
�
�uF���'�$��n��A缢zE$T���������f�\C|���P�Θ��#��RY��819���I�<���o��C�XǼAZh��+���Lq��M#,�X�8N� �4p&N}}������-�m��c��+X{A�������>�=�F-����kLh3��X!�����m{�p�{jf���c�����y�BE�f�#E\L�L����+K-Ǝ,< {n�0�Cz;��\y�L����M��2�����:����Ck��}N����������TmJ��h����u�W6���߻܈���1��E{qa��X�z�*35�	 � ��C���}��E�jʜ7�z�LhC"���kGN?�x�&'��+�C��ܷq�/`���
�������y�J�W�@��EB�_�#�&S�����?����
�1F����ӉK����"�&8�S�[uB�b
�T�2C]+�I��ty����,��@�x,@̺��7.5v�/��>* �/%.�>�V�^w�J�#�x)�����S%[|�/��;�o~� ?.�,��&>|�l3��t���Y��������w*�=E���� #��sI�ƽ��FD)9�k�B:���IS�ݻB�]C�W6��;�_����x��r��y+�I�0���ɩ���o���|Ȑ�F�]��
գp,��Yn�u2r�ע�à����K����z��R�,�tEҾ)����{��؍���6�X� �G�G1um%$L��I�j����e�0�X[Kv~�>��w:p�z���ar���p=�L2:��ݶ�풏X�d�q���]�#*\.�#�ݪ�+_+�2�30�r�j�������<G.�~���
oBյ�]+Ei�׶2:�z�!y�P�����k��]���t�A�TI�����\)o�{@\�F~����2��_�k�^%��(v�_�n|�-O���H�Mhs�z��Iv��}q�k ���mÞ�	�]���@�؛����,�w�Q�qKaa��X*�R��<:�J�S�`�W�iK���B	�C9�,��������D��'� h�o�TI!/X���M���5z�ڷ�/�Y�qĕ��\�C^�����������ג��$S�ʹ3ل#V��r�O�ؖ�p�w�f�t��}W��S�\�+�7\�N5���f�]�p�"[T�D��ۏ�_��uvv�f������_�.���{�a���W����>�5�"�KZ~���J��\S����^�zspГtGW�� 7;�#xq��7XM� �i��D�F��u+�{��|����[����{��Pp��J�����Z�?��=���4)���a�hz��GD	?ݺP��	-�VO/d*wM@M����
<fBU����eW�IYɺC�1u��S��������5���H�X2y�5V�@޾�+�. l�5�aeƄ[n5aM4�Ɠo���S�q����|�ˉ
�(Ș�����K�Ԉ��� ���/�	�v�+bkF�Q��#?*�Ԟ��vШ�~��|�����xA��R�~�T�^/oQ�0e�����Ƹ��������\�91��A�No��?�bR?]Į��)&&�%���e�U��ѽ��3�2���$�}1�DQ���[��6Å3!	9�o�6�?x�T��G��e`�Y�-+,999_�\G�͕"��.���܁\ȷ�X���\���Jy������Gp��L_;��y88�䎳 n�����*K[��+/S�_���3n�)�K��H�[���?r���u�#���<V�k��s���2�(����B�Vl4U��dqa�3�
f��ʄ�X�$;�',�����yxr�RdY�54�D�>����ׄ����O4ϑ�m�G��"��ɗ���P��}C�Q��sؔ¹
l����A��'ob�pw�>A�q�7��{�8
�hi���8A���=�d���~���$�Y6̄Y���e�^0g��}�-�˸R�ޑ��m	���8g�4�ח�ó�h�3������>7��>�o�9CS��5T�j繐G�B��\�3ԝ�����`�}M�e#�.�vK���*�]�������u8>F������e]ԿC��u�O�L4�.��H�*�nޠE{�F�uӏ�E2W�
/�+X�	R]��K�)�B���W����u�?����7�ӝqoI<��v{�e+�'�x�VU��{�h����=��:�eQWV��R�bg��vѾ�Uh'�n-\�Q�/m�
���&]f*P����8.(�����d��:3��	!��â�;����7X��>r�~Tu�=gb�Z-�>_�["H�n/�a���K�{<`��,:o�;��ci�V`�,�h*�i�XU�g���^�T�bsr(V�D�����U�_p���K��ÂABe����f�:���q�?�V@��RQ�L`na�ix@�Z��ܞ�����g���.Kp����Eb����]+kd�vz�����,�>�;�I����p,��Ç���]k%��$Q}}}���:�5��9�E�������r���Q�t-{䉵d��x0���>x�<K��3v�����0��m�� �����y��䃔��&뢗�'�����i~F9!�UH	4�Cu�1�� g�濖�L��؁��Xy�r�\a�V�Llnn���t��S�N�-l���'hӷ
�� �;���/����!����_�	N
F�zf�����dt�cFA5���^�UfA�Zu�9)i�lA�d���WTo�	z$ ��F��P���n��|�����B`�N����G�Xg�dLyy"�>�wB��߇��\PX�)z���2kH�E��Ӧ�;��#�:���t}�6����5��Kd�����}��X�L`��.��~��P��&=NPY�N�n�,��/�|���S/��g�/ʮ�vyX���]{b�滆��3T�d=<�$�Xr?��CF����gryX�ԙ��i�����*��0��e��\;"�ps;j�jr}Hr��%�6����x�P@����i��=�]��pK[��[J2�R> 0�7�BKl�/��/
�K_��	��t��C�LNNc�c���q��=Q�󆼞��^0��Oy��Vg������ e�^,N�����d����.+j/h�Nq�6�U�&���Z�fbr���`�>�&��lsFe9�X����[����5)����Q#�|h̢+� z=i���3.Z�<11QǔȨ?�4�� me�p�IS��
S���Y ��".`��ԙ��\��ҏv��_l\\���n<;P�Ԕ-�Mt٠S��(�������շ���`N͆�_������q#F%4?�:UFU������rz�]���~��\�[M�n�g���>`�S[[[��;�����Ph�67w��7�39�-���
���CX�3��yh�R��j��H�tvvf�'��X4�<`Jj����H�?�+F����^;pr�����e�I�+<]+ �	�zzzZh�t�B]���@�%SiQY`ٲN�\��R&'ݔ?h����:]�V� mu٢�f�&sh)�fK{�=<��P��-ҐM���N�@�~s�5����qxju�K��h��lv�2L�Y�ͨC���{�3��
9��S ��(�7���_�+oI%�b**-�X��(ⶵ٩I�#\e��d��u�(]PQQ���KNO�+@00�Ծd��|�UN��DGGG��V��.�����)���n�,Z��e�nL|�tG�e��fuH�����8���>`)\�کEq�F�E?�����Ō��f��i��"_���(5��׆<M�u��b�B3���<�C�j}�x���އM,��:r/YF�\"��"E���=�v����|b����R�=�W�ta�޶�璋7z[��~�y�Zٛ=H�^�C�o��)��s���=3]���_w$�;o2p�8������wށ8����GyR;@���v�ꏷ�99�������/�Uȳ��>������y222+3]=��'`���*�����CCC��&�}��:wy�?���9���������_h��K��P6��&ݴ��ٓ��̃��%c{�K"4�Z���4�~	B&���1rUN�h�td�#�GPs�MH�3�%�Lm�jӛcb ��q�t�����c��;��]�WٵJDPWV�+��.J=Ӆ?Z��N�3; �#��!��1N��iN+�TZ@����B�vu�-7������k����p�?�꯯�N��y���V���o�w����bS:7��Im�����M��D�����a�����_OA?*�<;��>�f�_��'?I�x;9�Ư��S�c�Ϝ�{7E����W\��h�	xv��ġ]��rq)Ĥ�9��t�`3G"E��$�����S�!�>�D	�%�B��|]sՇ�<����K���"���k���p1���� ��vK.v~�D���G�OS�ͪ��瑧��9�iԖ�Vw�,,縕Y���r������!o<_	õ<����+��������n�D��7�_#���NC��V��i��|�n�m��˜�6q�&����P���Ē�.�B9�����΋@7�!T}��ƊCW��Z8�۰�&F��b���\���e/�;���0a�6&$�"]\\ ��(,\H�K2Щ=K4��w%����&�%ʆ�25I.�;��U���#=�VB��°�F�^�ТT�"$�z:�5�:$N�8۝�a.��i�n�C�u��!��5���bJdVݥU%R[���s-���}��\6�	��!�����՟�yR��?_5��r'�"W����=�:İ��򻰨�/[��g��ot3�55R|!����4%u����r�����`sV�>�p'�Oۀ��M�ŵ�!"�8w\1`�<�*������g��W#�^(�k*T������}q�%��w*����*ɸ�[�Vi"J����ݔ�aQ��0Y���ɧ�a�E]��Ο���	I7�:�����ܣ�G�(�[_6Z����X�{j��y˗�g�Z�U��cw�:�1�%VI�G4:�p�
�vy���ĕ
+;��0i�_��Z����6�M�ǒ�
/�<��@;�DݶBM�U_ Z��՚Ҳ]�>�2�amu=!;��1�g����/5'�ͅ��"=�s�k���v*���G�c����9�<��?��O��s�d���m-���}zG�e��02R�R��}�*��_��5q4y5aC���G4��R����e���W̌����������#oF0����~��Y��@�~�P�vrPk�V�q����|
ћCB�~Jh��GO�r��-u�PIԅ��K����ِv�Z<�ʚZ��M��8E��v'^�48�@���JXc�	�<2"d+�c�����ҹ�4�$�{W��z���>}hY��R%��5��~�q�h�Q���k.�y5
��wv�W�g����ɗ�%+]"X����.��MW���R��3vp��t��ދ���T1x5Z�h�n]u>D4�צJ�ۇΎ+*T��\9���}���i����|�|����(^���s#Z�5�]�vэ���ĵT�Q��]���-�JL�/u|q��dKn�bΌ=Ito�j�S/k���E�^Ws�:�)������UEBN<��R��z}�å)�҅��i�7�U��o�opq�q��e��=9�NC���mP��o�󸈫0#׮È�O� �y��+�ֱ�/SF9���c}!ޯMרH�`�բ
9g���(�Ό������K�M�|q��w� Vr��$����8i��ܝ�;��W��!���@#~^���
ǖ_2Y�C�7H��d���uk�B��X��,ת��{�l�K�W)k�mPͧl%��bdi����ң�LPDs/GӪ�t�m���m����XH�v]�&����wS��?7, �=�Y�пw�/��W'°K�J>V��>t���O�	Q	��+��oP��l�Ǘʩ.�f^�(_ݒ��͂۴���9�}	��{�*��1ۧ$�g"���XW����Cj���9*T1a�T�]sv(	g��R�¼h��-\�yA~</GfKO\N�y��O�0����%�cɆ0�A���Z�����G|��4 �Q�W���q�������=y��e�zf�I�\L^jG��\B�Y( /�{�J�w,���	o�'���t��g��j�M��MT���m'g*Qs�6>��"�ǈ�xo��:����sTH�W�l$�{P9w�[�U�Mc6�of�Q�𴮾�Qu������_0c��+�/V�����[�9���l��G��5z*nI4ή���l�<?3��5'��:�n���&�B*��e)�	}�#���Zm��WI^i�a��-�+�o��U.仰�u~�;?ZC���Ĥ��l�
�D��#L`{�s�7Ҫ�b�}(�4^k �l�'[�l��\h��$-Qo2��T6��oe�����+����z�������@X��-�8�]�i�\z��`x�3^#�]Oh�u��Ls�r��X����V�#�w���׈�\]e�H8��QMu�c55dlQ�㫧��)�V�p��2k���X_���xZ�o#n�M�Br%�$�ƭj�V�/���r���N��&�^���mw��*/����M�x�c�cx���������7ڙ���.9������a�k�H�å9/�#p�7&ν�c������h�	o��PO��S!�҇Mn1�B�8W�RH���K>�_�Q�=�׍��Z;#���g%�G��l^)V,����-��yiɳ`N���Bn!G}���15/qCy=&���4�����dM������	�{R�f��Mѫ|���u�t �`���OA�9�wh�P��8.�g��{��h͗���Xʩ~(9��*�u`I�r	YTekd�qA�4Ds����ͬ���	�=�nհ���� 7�{���BU��B�����w|�gA�:��D�l#��t��CIw��ê#����β��Ȋ�e��RM���v�q�gc��c4�3s��^��b���h��n\X�@�5&��F�/�5�����S���ޭ��f������=xr��[���w�i�8��61�����!��6�%'_�kظ9	kT���;���plX8F?Y���9��Ԫ���P���)1{��� ^�YSs�B���2>Y�󎭭�y)-P瑘�m�vcU�c��G�x�����<�q���޺T�5I���Q1N������;����k"q�.#�zzzK"���YQtC7�4ٜsaxm�X��Ƌ�J*��|0Io�F+WԻ���z4_b\�����FH��f��������@1��:��j$Y�.��+�!+���c��ѹ7A��!5,AK_]�\�_1�0!�Zc�q
1X[�#�&�sL�^`Z���)kw�E�W&ʀ�WY��h����,����%����j$�ZV��x�$Er1����.���[#ۄ|�(��p�Y%a��Z��DZ�g,`�q�ڧ��.���^t#�m��'\�4�<�e�
4�<ahZr�
ȝzz�]9�)S,c�(F������H�<�-9hX�aA��#��lT���oe:Z ���9)o��f
X��լ��W9y�^=w!����%�O��G-��8L�����ۡ���-�p_�3HC�� �)5v���9�CV�+ҽ[�������2�S�u�QUz=�x^R�Sc�O�	C��u��~@$�ߕ9���<�?�R�1�	4�d����8x>�Cn�xn��l�xt�7�X�#ӷ���Q�Iŷ�ͨ~mw�ʍ;��ӡe� ����_�8C,���$�4(�V'2�8�hiZ�ϔ��� ����]�Xl���[4j�>��]�hğ�,'Ʒ���3E�+X��ي��uu��k%���T�;*�%��#T6A��NC�߰��kZX��\j���NL0��`r���Ṃ��'�@�d�����\�Z��r�v��%o��s6�g=���K�$,�ñ oБ��cG���[�l�<�#x�y\�(��[��j�YR�b������m�@B֭釋0�z�e�j����ܱ������)�f���c-�<l,Fs$b��7����69)�	�ל�3�7�1�T`��]�.{_h>yQG�2���Y��y��.��쒳��#�|/K�]�cā<����y��
y�~�4i(�@bg7�rYG��N�r�զ�e�<��E^�䜈J�=6��E�o&b���C�[_���l�a+��?+��d���v)�r��k� a9=�Q�
t$"��	y���5�g'�ȘU�ѵ���0.����f�eǎ����o'?C1�.j�o�
T�4켒e�� \����3ɍ��4ߚۯ0�����=�Z~�ϣ�J�0���A�E��Z,�F[�P�AU�؁��*;�P[�Tp�����٭C���)��������Kx�\�ĭ��܋\L��9��ҷ��{�Q\�ّ8��;�Y��<��T+�a�ǛҷP����I5`��������A���v��کk/��o_��Ӹ݃�|T�(ˋ�.�'���ߏO�\#�����{���/!�`��{�a=I���KA��r5]"��.�FJƥ����B~���U��Zv�Z»�\�8w ���U���9<h���c��ނ�ԓlmF����	Une�������W�@!�kڂ_h ي�ra���03/��w�����{��U� D��rg9�D�~2x%��������@<��T.�g�%�/L����4�`��S_-��^.T���ު �9b�8��� �����tՙ�z|�A��*r�4u�7g�Z�36�7Ns�]f/KK�X����2i�o �xy�d��0[���Q�����L$Y�JG+i��EP��9t=���r�k,޻�2'�9݋9�W]ϧ�`��F�e�/�:a��z�a��Y��w��5#��6���O��X|6��=���θ
�@��Rt�W6р ��Pէ���٘-f�����bV��Ǐ��ܤ��
�ζȖh��I%��#����*�PY��6����X$%�{��,����R��C��`zV�G�b�:�1X}۞�~5�4)XSs�]~� �|��k6D��,��R�Hҡ΄Zua�@�D��amHUE�9��?��A:�*�hQF����^�a�����@X��_f�z7a�k����ـ����d��D �#�h+��0;+y�tLP��֜��������0���.�w����m�m��}@�>���ʒ�wu�Z1����.�[�W(�l<���?39��R�j�{���Jl�����m��׉�%BCbZ�AM����D��bS�*�u�z�V�q�5MBoRԕ�,{i}ix���İ���~��'┋Ͼ��<���k }�j�Y��WGA7�݋mN��?�M�B���[Z5!�4��^���9���`ԣt3������0�z���a@��P\��bsG�����ʂ�k��H��<٢����`xu���|�Q�R�՞Ae<=3R�&�l�G���}Z�j�M	��d�@�"��Ճ�CE��#��4ݮYH�K�T��zh�[�J����(�p���7R����*��m� ��17M�Z�H�2am�O�����1bq�$mc:G�Ve�sd��."L�G$UWc�5��4��!lY�Ӆx|)� )-�<|��ǝ3"Q���C��[��Lu�B7�6��a5��Nꌊ��J���a�4�3�uQ��bQ�yM�e�����f�95u+�x�����h[Ȝ��㒪��5ԵӶ[�Z'������L� 4)j�w��T�J`������1�2£��uO��Uq�-T���Пcgq�;LR^FA]P�ܝ�Ea���[7��_L̟\hԲ?_m��c��EGPO��)�h/�*?�GF=��6 �ҡ��ߪg�y''?��]6��ز��73���*"�����1+_O�(���^�i逭���/�h-)7�(+�����+;PR�.���Ц�����7m�^~���q�7y�j��X��G��!����?��M��vJ�4���wu4��C�j��2� ��>t��7Q^@Yʻ�ӡi|��v;��>J��u�OQ3��5sV�Z [��j���P(����
br��ۮ_`��vKX�C.�Dc�gC@r$�IK���܊��D i�ޏl��>�@u��"i�/`�k�qg�d2��n�G�j�5�(vv����C,P����Q�@�5��	F�7�k��Ҩ�v�A�?X�vg���/�U� -_Mwܑ�7��op�����@��u��	M�.���<�ܫ���5�)���F�NL	 	�(�F˂�2�q�G�W�4����0F'48���H�`5��V��YTl��[���Tax!Ǥ�)�����R��(���?RQ`�>�q�`�a纼��]��.�՚�p

��J����l�����+��/\�Ҿ����L��Wy��H��Z�R�������J��ƨ������v�+�[8U�V�Q��)/!=�5ש��N��;ŧ���zm.�L�oB�Ӊ+�f�����A�l�,��3�i��ã#��WR�>I�3 ���9�$�h͈��O��j��VZhC����^~U���U����ZH�R�3曄'V:�iW��}&�Y��Y�^,�,��ʓw��
l�L����G,�l�	�1bN��&X���kX.�?$x�@b�%P%]�TO1�����P�ˢM�k!���[�^|�;<�I�h�>p��͛�;�U�RKv6�ޗMO��yj���%�K�.cP��k���
���X��]u@P%���c��`�P�%^ JH_�N/�f%�i�q��Q��,O�q������+Xь7�/}��3A���iɕGF�}F����S��u��rer�$y05E���kt�'MF0���l�F�N�v�p5�l���.0��:֬�S�霐�ˍbz[��bH�E|�^	�c]�,P�3����6:��R�ԟ&=��ZF�5UC<�֯_��6�Ar>}u�-��1Jڇ|�㿖�k�Ԣ��ÏT[}��&����4�&��yR�;}ݨ��*�Z[�e�!<i�+P�P��^*Zhw�.����[�f�M�識�1A��r���O���T�r8Y}�ՏP
k`�@.��q��z�U��(f�'�/y��<�_���N E @i����J�אռ����K��H0�m��x�����5#t6�L�
V�淐����8Uc
�8/�	X�.1��h�%4�Eh���v=����g��2�6�Թ�q��=L��j�FOC��4��N�Gծ@I@�@`@]ZI�@g�ݾ�.�R�F!շ��V�=!�#@�^tC�����ٍM:����By��$�O��(4h�n�"F�M��N�M���lm�[E��z�:��%��}Y/��ش���9���R�H���gh�!�t�w��8�D�fc�w�q�hrv}���8�Tt�q��>��V�S�>S+�k�	�Mvx�7֥`�Ɉቘ������Q��U(�!�I6[��]��c5��_�ʷj��j��+-�ǫ��9�.>�幒��s�0�YB�JU/�K<�ڄ^{{����(���Z���4����P�M��\�`6�OU�R#�.�+����©�c�%WS����,K	�m�C���L��U+*	4�O�Z?�|�8��_w�
��+��\aD�I	A��������ܒ��|u�E~?-�Z�Bu�6�A\������H �/#s �W�ďjjO�x�vO��k��7���4�	���C��ayD�6���Y�d�����'Y9���q'p��z��B�i~���S�g�33�x�T��%���{'�!j� �O
��9�4�l�B���Q��V�w0�`���Y��eM��٨g����Қ�Q��'������^g����Åѣj��K�=��j�#HS�����"�!�+�;�N�`W�U���Ĉ��D'���-�r	@�ԓD��gG�B�\yWԳ�t\����s��~cE���'*3!ސ��4�pѤG1�8u�^���P���!��e�e�k�a�9���þ��l�~.Б��zFZ��T]i��+��τ�|�
�R�I2alY�_�'��?$1 dI�92n|VVǨ��-W�L�p�TT�)<��xT���]�bƆ.�B�JHN)We���{�%򬩥�i>^П�E�a_�Ɖ,�Bi`%��ƨ��U^}S���oT_�{��7�J���-Z3��{}�CYAt~!|��Ja��`y�`�R`�S��]3s�$�(��֯_>�6
!Tױ5aa��1�4ػ'g� �t�_̛�=�����v�u����v����gl@����1��*����ꗆ�M��0�[-�lxA;\���`ݼ����1�|p:H�]5��y���yŚ`��GkLô�a���O��m�k����13JқC�Z0G��RG��e��������D%Y� �77���gxAmWk�!���/����g�s�b��8W�|FY��7�%b���
����X%u��>,�֍�_&:�7R$��zt񵒊
g|�u�=䒾/=G���������Wm	��=�ԾR���RB/%;�d$�r��s��JO,���澄��ڥ������;F�`v�������/t�j��+�a����{���_\������_�����g������V�Ż�7PK   �|�X��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   {�X ���s� �� /   images/305f7d3b-a649-4bb0-9743-3edf8bc04acb.png��csfMۅ�ؚL�m��Ęضm'WlOl۶��m�zs?������zwUW��{�u�3\^N   HJ�(  �  h64����|Y�� c'��  ���$Q#�  __�"��n��0��j�d�9��ʁ�F��V�#u7�5�ƣn��50��n�?�cm$�?���.��=~����t��&a�̀����3x��e#d���I��H��+j��ʼ�W���\������U�|Y����1J���0j<K��=���&�9�7����<��K�QA��-B!�[d��p�+e�c�n����뀿��T��!?d�� *8�[����_q?��LPW��'���Yx�w`W��X��ꈴw~��E��m6�Q��V�ņ�Wߌ�m����x(≥��\�Q3����ʻ�ӌ��f�p	v�AU�rn���ŷ�%�1�)���'��%a�sO��U���rӶӹ�p��"��w�ʽױ�{xj�㋼4�(��4���n��c�7eu�P�K��p���hv��{�Z�����q'���20}�_gk�3�F'9_����.*[G�6��j)IH9�X|nR�:�?��0!�@��G���B��i��M�R '	3���Elh�X]	�qӢ�����+����&jqy(>��=���������Ų�1"�����1�~��%�]0���N5>,�Oǩ�K�\���`n �2���P����b��m��[8��X�3��f&8����4]���UH<��xa+������0Ӈ�5e�e�B��Is��>�����AT���W�mK\��}=C��ie�)�>��ee+aM|�i�K=`���OrƵ���O>*$:9ݭ8����)!l��g�S`�:U��j�,�균����o/<KNj܊�}����t��� x[�nɤ�Zr�[a�}{�b�q'(��W���O0z�n�0��� ����tᗵ�B��
4ɑx\�^9"��:}�_��IH:)��۽B�{o:sN��u��XZ:o<��4����׾��I�0�M0���B|�k�y���0��p�<����X?|�g��T����&��9k��}�lb�F����d�t��2�;T��v��C���`U�:�8w[-#O%>��N![��}5O)�e۪�-'f��4*=���ƺ�~O<���X�����(�1T 4p͏���2v�*�icd�x�S�����U���|��k��z���K,�Z�4����q���_�Jqk�������6=��c��{�
=\D�fƃ��p;�u���e<D�$���7��\E� U�6�ll��-l{Y���DG���ц���@�Q�%�o��z�hNOd OlVw\��W*��B��NF�A�~��qv��h�����ĺ�px��L}n^r�>��RC.�֏���l>|�!lZsI?J�rn2||s�jlo:?j|� ��g��2%_��v�|li$(�7�J�\�6���6��z��~�|��n�9��W{_X�J��9����;k����,�Y꼚i�;�؈����s�&5�O��=��L)2dx��ϑv�Kk��+�>!��d��W��?r+����
��L`gQa:a�� SYֵ����b&m�D�0L���V'\D� 7�T|T
����J/����%�'v�xڅQ�G�I��d�"]����}4��}�c�}��X�Ք��(��]�E^�D]��f�V�|a�충g�#��^��F��m�mg��1����Y�G�����}���ږ������˴�'�c7��c�9Ρ��H�����^ T�q�����
�h}�݄ł�j�ȅ�TiT`M�U��&Z��r�;e�1�*��{�^@j�#% �ψ'�$wcT�l�)9,߻��L�'�"i�K�D �Om��ǝ�j�l���r��`��[ru˰|���g����\�Q�y��cQ*
�3�_��V}u�Y������-"��4���������J�h4bb�r������f�-S��e��&�46hW<��u_g�����M!�E5�c)�T�t����NOx.��1�YL��������܂�� ��V(0�6F�
�K�n�Ov/�X�cPCP�rrb�u���[��l����1H;nE?#a��s��*��������q��ULQ-s'������y����rСsr>�B#�uUK��i�}~ֈ�?N�B��πgN�u?dd-"�%���̥��[A6%W	C�	�����Cm�	�/��Ⓨ�Z���5v��#��9�v�7_��&0�i�2b�bNP1��M<`�v%��>�!4~��9|�'�n�p?���T�$k�~�/�Q�L��v���G�� �VK�����e��*�c�S&ډf�Q�F���.��iZ	[������+#���Fn7���|����.��w�^7��ziM@-G�W=�'���D�?�& ,�uMu	�q�v��>}L�|���6\�>z�|��=�Z��݊�����n�?w������m���3�Uv��)3\	���t�՞��Ѥ���d��N$!#��TvO�9�JP����F��E�G��w��V >�!7����y&п똌Ҝ� 1u�v���EDm]qL2Z����揾���3|V�U�m�Ax�ɡZ�<�%�<�R��d۾�b�p���W����*[�4u�S@����Ll;!"H;/��.d���b m���ֽ-*؋��W|9<�cL���A����H�p�v��Qkc��[�t�����4a�n�_.�6k4Ń�6NZ�����w�Ӏ�j�I*��]YD�G ܓȗ�	LO3Z13i�oJA��-�����MX~?7b�aW�u��i:���.��<ls���U����y4���'���B�vy�n��������7�P�bP�3W�}�[�K�-
3G��z�Q���V=��|56-Ż5:�I%D����1�I��Oc;���4����!Մ��a��XBWW��(ˠ�I|�siq��gkcc\KK�R5avV�T����i1B�T�PЎ�Bs���z��ζ����Tp� ��J�|�PK��J�gX1��h'V͞A+	t�u���W�k�ழ~����I�,��%K5��ړ�F�+���U�+���\{٧Y��p�O�����	�F{5⎊sv�gG���э�&�~7���|5zle�k�g$M(�{J��YRu�	F0�d��`5�*n-�.��:]�dY�K�X�`�U�?�B�E�����<��yV�h�U���X���XM�e��dI��rz�����O<$�rjk!���Wi0�1@cu�]*+t�u�x�d8?���؁�Mõ�z�U��w��{1�t�]�؀vC�o���kʒޖY��ԓKOSk��[떸�ʴ�M��$�PH�B��SI��/�<?�޲��w�ƀ����6[�_U�]qk8	���P�wq��k�[��½�Sv7z�Ǟҍ��q��Qp��$���g�d����Y��3u��鱦�4�T��gDY�����nL��cy�Ƥi�C�U��]���2r���1TeeM���G�pz�^i�%o����3ꅣ
��@"�|L�W���E�Q'�f�N����81qpp�}�=u�Y�>�����gq��w]u�d�v�z~}~xs�O�0vi�S��vd�/��xv>mjv��|O[7�̪�!��wE1f�Ē����ڱ<�����*
��+�A�sA�յ����R��Q8��d3!���s?�21"FE,���1����H��FbV�+T�~5��(�^Ey���ў�33B�Js��Єܿ5lR����gw�;N�A�$M0<x���
��4-��Q����Kͦ�ߝ+U���&�m���&R� 3�Ӕ�2�-�.�����W��f���$�"Y������"��݁� =�;��I>�}(F ~�!+$$�c���ʴ�j���u��q��j�p(,//�,oM����oʖ����ߌK��lq�!��"U8��E�C�n�~�B�i,5�z�C��X��m�^��럣`LP���_�%�/��9|ԡ:�v�U�?8qp��BkW���\��e�����>n[Z��5'��S����Ҥ[����.���rqݴ��S��m�?�N�Z-V��:��5`ٓ/�,oA��4���wƨVW:U4����cFk�"ۏ�C1n��y��e�h��Y����t���hs��OEL�����ZRjA)��cӰ�����~�uf$}�[8�T�m��P��>9?g���I {؅F��dm�a�c�4�N[���+�%�|dB��L� �͑u�9f�֝�����Vtr��ӓϣ��4ԁ���o����i)�U��3��*�Z�z�3����U�dǴ	9>4d9֑?�o�L%�ڎ(Z���ɺ����W,�\��Έ�_L��g��/��4�&_�7��ӌ�܀�β�@�a7#+������5�9���7\]]�{���:��|�u���|?_�����^��d֢m�kvޖ�]7���{�|j��<Jx���Q�q�^&���XV�RљH'�)IOCԣm�GdQwE����4�Х`���l�5���s?��2�q��$��w~���5��Xż)~��m�!u8��/$�TFu�qx�o �3�U*D1�jPf�#��Q�"K�<u�߀�q�� �>̮�;�c�u���B�.�4-S�萍
'���ς�c�qvj�vm�aw=��Udnԓ�̈́3)c�D��ڛ�xa�Yq�ŷ��,��n�>u��2ʸ5;IL4�L4�j�9�(-�x^X�l�w�LFDMO���e��&d�6���,�����}J�G�>t�:0jy<���iW��^��pMN�}D�5��S��6r��s�;:�����3i���k#CˉM=��2j�����	��Efv�j�<鸍�O����wX�V/�z��X� �� ʹ��Ҟ�S;�l�.CG^~�m!J�O�V�^��!z���&���H �u�Oz��Z��o�����0�^$�#)�:A�;$����Y��0���8�r��<)���iM�r�S���Ӥ��2}��.x��������
��K�e?���'��Ξ}83^��xz�mga�vj?�F �i�m���o\li+�}�a��^?q�c�uы��>��c| زj��=a<c��T�[���e#1�O���V�X�75gP��b���� �8=;�T	C����f`��;E�S��.�����r.�2N_�6�_�C�_�
�`!}������xR��H�ӂL��gT�b��>.�h���{b�Z��&R1�t�|lso� �?��>��C7*Z�O�p�	.G����a���#L�F��Go˚�:�Y(s�kxXvx]���]����ܦ�!Y~|���{�Xk�YF<�V-�J�*ǉ%&6�i��������mN�'ot�?��5�т��Ƈ��,�^�^�����ٔcImQ�Ah���Qm��0'������Lo!����E����/E}��v�z52%��RS~���g���"G/�j<*<�L#.��䤓���䝴{mja��o�O�n�l5�,ЛB˰�@\i0O��I������h�c x��)��$��\����?���I�vqro�C8�Ä�c�Nf�\��TS�|e�UC��.7�|+|�5
���3E�5�H�I%�"9�N2�j6�zX�lZ}�<�j2m�S�F�����6��'����uT���I�ک�ge��(��1lC��M#C��JN���e�f�_�OJ&���{�韔�Ih���Vc�y��i�ꔀ����I��J=���n�]���ݮ��g�6�Qna}��k��<&����s�د�h�@�Ql���ʼj�9ʍ;I����z;�K�r��F'���;V��,�#�����2��ˎ� �CiA�6D)؟f��FZ���	��'�V����q��\\a�E�9�&T8�_j&�B�����6�^����Q%s�-����e�F�ލH�G���O}�9U3��c���-��չ��`2�<d^�F �L�j���*U>��Y9��� ;�l�8~p�-�^o����F>~3���|8%ι��WW��ҫX�t���%� M��!���J�AZ�(�����0�_sCݩ#��T.QȦ f?�OcUA���Hw+�ι�W����*M��Ad�K���jH~+�aQ�G9f���!��N����D�`���e�Y��|��%�Q�d��
n�>\Y
�J�AY|���]�п�U�_��G����m���kX,���!�{�����&_��@�$�Μ0l�њ��eSS�c�GN���.��!e�~���c�����:��{Q�"��G���V����w�M[���uk:������!�NV>O!k��O�4B)�?���߲?����%�@Jg�����fU�62��(QT�\;�r%���MЉ�P�28[(���-P��S�;����Ȩ��L}i�Y^S�	Ɔ�J$[I�V����+1`�^|� ���L�Lؤ󹬓ެ�	W�?c��g�Oy��Zm¶Nߪ;��wB�BР�����/�Q?΃�J14�5h�~sA���X�
��e��Ƭ{�VT���9����\ƫ#�v�r����_�h�a�7���i�J�ƎE���FU�-�L)�9�
k/�Ǫ�.>�U{�y�� �ޞ� �o>$�����d����P��5K�1g��2ef ��NjE=�
.�5�MIi��ۃ������)��{�CM$;d�}r�@�w���xi�ʂY3�A����@*�#E�"W�&�b5�y��D�f|R�>m��I*{�b\<�]U�*%�VR��bV�g��_x�]k�"�@���@5�� U�q6!+�%	ۧ/,=�D�|�%���z\!_'^4Q�j�>�c%\(����.=�ǡ10�n[ˁss�Oo+�X��f�$hƤ�������U��5��|��M�V7ý�	�p#R?�ߕ���t'!i���p
���u�?G��S���j��S�B�q�zd@�����f[��a�HQb���_C3��'2�����+X���ze�����'$XiK���ďf�a��z-��}&]��ύ��P���~Wb��̓�hT�q�J7#�?'ޒ�'U�x�4lپ�$ʁZ0���<{1Z�z�s~p/o�z���NL!��6��q�\����E�����2 �n|3\d��d��O&��]|�A��Iqο�b��^�u<���"��?f+�h�c0�=Z��]B������9��ٱɎͶ�h�\k�*��?��Kg]~<��w��-�p��~�郘�C���.mêyq'��� �矒~-��<7��#q0���I���*]�a2�����$����T�M��Ha�H}��Ր�WjvL���p15�Ux
���&M~G�칇��Q�(]Q��I(�˴�_y}�[.7�]�D��|�,'�� ��+�}? ���S��=��n��|�L������s4��)�**�����7����ͤvv�����8��f�.��gF�%Nh�,<뤠�%H�J�rH�$d�
�V}��M�+gn����ϣe�ӇW�C�� ��[c���	x'��)�˨\i�հ�=���!M$I.iI���qu��͢����:?B�ͫ�����nt� �ԟ<)��֓�	��(~��.ڿ�^���|ޒL�tmJ��xz�� ^E�� ����zez3!�Sgu�¦4J��Uc��y������cvF��/�_�o|O�kF����)���;��m+9R�I^�Y�Ύ�����~��Q勧�6m'EH����0ޗ���%ن gJ?����<��|���oN2�׭1���cSΥ>fAU�Ϝ��->K�Җ�l��s�~����4�zc�]����o����5������6�Nwqc��a����6�f.P o�E���v�K����{�f�`���*�ϣ7e����Dg��t�]Z�x����ChY�gc�ᶝg��	P+H��p�d�0_��f�ع�k-�H�oŗ_�_�:ʨ���]]��c
Ά���̭d�K�̂(����W�I�d	��*-���W�M¸�޳{�ۊ�3M4j�y
����y�.���\��l��k�i�W�����A��q�BAh芓���.�fq࠰�5�^���0>�F=��5��W���{���ش"s�$*�τ�"�����T�����d8��!������:kW���}��y����ޟ�2�� ,�Ap�[iu4��G`�h�pɨӮ1(!��ф���(�e[��Jx:�H9��Z�U�on����Q��u#O�Y5}���Y�������O|���\xi�2�V�/m�sFg��J��0�8�x(ݾ˶�O��Z�2�oD⽟y��~\Q�}[]�<ݸ�y�8��$���NH?$l���P|�7��U19p���=��)�R��O.��Æ���)��:U���:̨N�g���s��w��!P�o[&Z�Y	V6� �uT6�ϖ�/�p�h"�D�b�q�6t|0ZoG�)H���@�6M�x5eUM�q~X�IrC�J&^���D'w<#q�KZ���1_�ԚMV��{C�3hH��Zޞ�t�>�l�&�x]7ݏL+@@-ɸәt���o���>����O8��PI�B�'	�l~�[ƛ�;6��L�1�,�'y�A�?w)�"���I˟ڑ����f���+Ձރܷ֝}�Ib{u���?��2{��"��7�|�uӡ/B��7������j�z�0����t���9��-�q�}�������i�L��t^^�?���r��zA�7�����&�{����A�RU�nTU%�h����Ϻ�£�Y��̆x{��_R�:!�}\��^�m�ao���ČM��v��<:������i�"�p��	�a��}��`���o�E$�$�T�r=�@�T[Od�ݴ�p/z�����:�1�roMR;Hj8&*���>�/ѹ�`�>��s�X������l����r�@Z�fռ�w9��铮�E=ѥ=�d��}��@U�F���W:5����#���t[���FJ��KKz�/V��}�T�҉PO[��	�A����9B��ղϩ0x�_0Sr����K��!��4Q�jeN���7U4�o��Y��p�a{=��X�AH����"����?�c�4�>�]90Be�͉S �/�-�x����v�eG��wm�f�w�%J4�⟭��Q$��k΍�P�r�CZ���c���L�m3�1�x��9��t��z/�V� �<�/E�3ly�c�F.�?8	b�}P+�B��M��J+R�
�4��6�=(����@�!%e��+ߴ��s��J@���DwIK��Z��0{Ja��[�,��迷��J�'Q��w��g3c�E�1������I+��ϳ%�7�\P��6q�K�ͫo$�R���^Pdi�*kPQ��l>&�c�CB�*�=���c^�J��5��P�\�
E|	����I�L��<��C$ ��!#�qQ+I�&J�C��4;:��,@��[�7"p+?����!�w{�w��<YV����Q[�@��r�	�Co�W�<�*y�ls�M͢�M%Va��
�~}�q��Љ``�7_}?�8h����'�C)�=R���&O�SۊϞ�	?��������2��2~L/ńT�Y�WΌ{�ɸ���eЉ�E\%q�BA���
,�/��3������K�C��*�fv!̛5r�!��D�/�#�QM�2QX��*3�۹���.����;���dP}_ߴ�M���=���@��_���s��}.�u�$MRdH��>A��ndn6���Q�.���)oF9�o8+���K�H2�Mށ/ވ��tL���ť4��W��q~Lf�E��-8i,�0c����
�2�y}� ��$h�d�Wa�����A��7�!9��jW��ڴ �S�g�L�;���05�{�-��X��#��b��+������ ��
�ԂYv@�q>!�3^�@�U�q(K�a��=�e�1r�&yGr��@�5�c6���p�(�
�ll�u�A��8١�[�?�ZA/6�>�5��Ť���f:E/p��RZ�bGe7���0
r���=~C*�-�^�`EH.񼹴T<��#,�"�p�R foR��a7ty�(�*���+Il�¹o�b��S��f�����l���0jا5��\�J�s2t��H�N�(�/�6�h'~�M��x�u�X�j��W���i7\D	h(�+Z5^����Q�rRE��:�p>q+����E\q��0f,��gG��9� &RP����I���p���{�(}�c�H��ˮ�-� P��H���*ж\";�;�[�(wb�S9�F谽"ݷ�A?�hx4��Ҵ���J~,tM�S����$�K
`�F�X�A���B���m��$M&��,�X��sa9!Ǽn�j		QL�ٓ����w��C2��);;;��{&=���2�﵋`�l�F��U�]�pI�!�f.6L�r'��'��Pۃ �%��)z�|"h`j���B5�����h�-�@����6#hF�G��ʄh�5��q�KL΢S2��1�U�Z�.Z��b����X/�2��a�i�M��^��8`��}Uk��Wg��jU#��#�P5k���p�+1�����h�oy5d珕Q��=��*�/��ZOȍ�wr�+�nD_w��-^C���X����r�ٓ�F���a�U���[^�d�0�E���k�n
�p�j�C���Z�Ժ_a�Z�4t��h6�8��6Yl��>7p�S*�p���G���k$3P&DݦT���z��]���Pe8�Z4�xF7�P'�h�`Zͦ�%�|�����T7���:�V�ˁ"%!  ��UHV 9X~���.����MGP$� ���0���B�b�U����8�)3�-��T�^��5j^\�$ݤC��d�T�v�s
I��`?a0�L��:�f�]�*U�j^��̼ ��㞚f�� �#�[��XE����O8Z.�Z��������!p5��+�%3.�Y���gn�����)�q�n��k>�x����/I�
����e�?����+���C-*�������~p~c?Z���
����-|,�Eü����X��7�v�`�t��6]�/��9V��f��܉�l���t�<T+��Ƌ��&Dɂ����ۋb�G�u�
�؎�hNy�:-->�r��9����װ��N�ςZ��	mJ|ޓ��DA~nmy�M�Mre�S[�o�#+���>���W�I�Y�p<������BK�={�cܯ��(��p��v��%0��c�-Ww��C�A�K��X����́�H���X�5ݤ8�<Hѭ��?]{�t���-�p��v�Ł��9��t�V�� �7�(���FlNFC�2�v�QQm�-�f&��ơ��"vJ�=O=�,�9{gx1igJ ���zƠ�)A7H����d��6�R8�����2b�D�
-�?��Q�3�~��&��g;�XΚ8~�a����(�8�Oc�7h��P�p �ˏ�.D`t9mV���V�� ����A�������F˃o6QՃ���	��t��@b�:~�~�CO�_���:Gz����Ď��������郣O���z��c�m��;��z[ ��n�@�B���sܔc���Y���s���JH^�Yy��l��!t���A���jh�j���JQ��vo��ISTR��_7�}�'g\Bu�y��
�fz�!ڪ�2�l1Tg%��wx �'�T�:  �K��'!�^��֌L���H-V�V�_�F�H	(fFtF����8e1D����6��#�&���<�ޥ/��.����X�-���m�l=�e->^n���i�v������f�_ h�����oAr�=�n��|^xK�J	�?XX<�aL�#�5`�(Ƿk��_��Oo�$���6� ��(� �Jź��U�YU�k=��<~�6I!�kvh=���ӥ\eDx$v���]o*/t����ol���.2���@��U�jm�d�!�ϛgվ�mk}���g���<�у ���q�v{�^#���[���3A���u�_|P��U7� (�m&A\J��5��u`+�..�^̕��S�Ӧg�%;*�4܍�:ձ��� Ȕ�8Kђk*ۿ�wD�bF����¼⠀1G/f��Ŵu
�6uU��)�^��+�+τH�5C������� �_l�4"�㸃�6�Q��V�	wqq�i݆�?];��{ +:t�ږJOo�t�ژ֞��>n3�_2^�zF���N@�U+��8��bV�*�A����d=�@�1��;�.̜��f�9Xd�{�*�:��H�Qg�	Az��6��%h@�?�.VB�$���C����1/I�S$�gf�=
Jr�y���ƞZC�n�\}��1ܓ�
��V�*]��m|V��i�.N�nTT��v�W��&@�ƙ��H� �U�P��Ȥ~�褠6O��km�P �Qm��گ����[�� �����l=ʆ�G�ձZe����b�%36��
u��N��{f,ʍxg$Jc+���+u�
Z�2�b�Z����Gǹ���7�)^ ���)�UG�,�_#V̧�5�ȴ
:U�]%DB�v@��`T��n���ǩM�u~�E���ώ!��ǰ���wؾ�@��{�8I����"�Σn�h��G{��8�O#X�,��&J�t��W�����y1�p	�Q�#��ːF?�6�9Ӈ��"�#D����8�Z�Q����]`��n�
/#f}0N����rب�h���R&�fP�$ ��T7��7[7|�:~�dl���)��T��_"�P�sVL|H	K��ٳzX&�0^���M��0�S_�ް櫧�D*��,��1�E���wj��̈́�>�e)<�I�@��B�����L6����wؑ+�љq	�
�2��mQ}/�7$��G�[0��^��~�kW�#�}8�� :�m� =$�߀>-�k�J!_S�#�h,���wh fL���1αx�lXG3������ҹRֹ�>�����u7G�E�e::���o���u���W/�����	��x���ۅыu�(M�TN��3E��q�qϾ��p��6\р���1�}H��*O_Z ��L�5�ڢ�\��ُy}zL��u�1��b�0�I�8;3��D��n��]}��~�7;HΔf���7�*�=U�W�]
����.���錸�d������g~FK��céը2͂�_Ũ��P߸
 (�!����0���>z�|���=��!�XC�k��f0^�ҳ�I�,���`�5�����[��C]�Ab7�L��'x�jYh�����-7�ӛ%r3�9[�!b�N8M�̫�ؒ���r�������i�Mv�.�Sa@z�!�Q*.V"�N���O�Ѩ��} >�gS�H�r>v�����IR�ӎp��q[W�J�R������UYNO�A+� %��eڱ�3@�1���W�Κ�����VJ��(-�����xD���U������ڃ��l��"N�Fb�_MՌ%v�줄fp9=ĺ��;ed9�l��X��}?!�:�p��0�HQ�� v^�K(e���ᇏ�������Ǎ-���x�96������T0�6v��a�&���j��a${�<�4ן��XK��8��+ȴ�܉4� ]�:��ѻ]���}D�z	[iIۂ���sYhUyY�|;fT�@*�Јѣ�օP�]t�M�'��u.(/\�E���A�/���7p�!�����Y�Z#�CM���ue$�b�X�63up=�b�i4��AY�5��|�9�p��6ēsj}6��z��U�,���;F���0Ǹ��C�9�����ioX�휯��E
˳ML�ï_0.�|�/�M�~���@�	��s��Kpd��"B_pk�j�=8" p�:-�$R�@oG@$�ʚ��U�q9��P�  ��~��hlr4do��R����0V��Q�넯��<�85��wl��`����Ɣ��.���7���s��%EG�ȵ�j�G-�><8��ǂ��ˀE��f�}Mx�}�  Yvj���l�t�4�㠸��}P�U�yk���W�G���E� ��y���Hn�׈����BZ���C�`"*���ϝ)iv�D��v(,]Vt�l�)�n�JQDjBwx��_���<�	#H�nWMQ�=w�}$�� ;�,mR����������w�Y<����,��1�*0J�J��H8P�Ը�Bc!�X�#Q�z�@�>}\�%zǟ�'&q&�t:P��q�*�7�ԠS�lV/3��-�%��.P�����C`��t&/4��i�8Q�P�u.e���u�l��q*8S��z�GY��F1�M���$�&�{�����׊~]�!��|��ou�DF�6�eд�����v��R�3{P�:R�����M;��#H���WXKW����x�1Jԉ< ��=���dm��C�2��U-�+����h=:��N��
'�LQ�/	�'-�~� s�ѣ�k��.�N������C-�����4ʞG+!�5گ��1E.�c�:*�"B��#%�4��=jQ��%�A��n�³�c��/������Xm�MPT�CD?Ȁ����A�k��ʑ���.1�"Q#�
�Y��[�.Ɩ�Ո@	�R��2D���R@9�Zy����F2�DA~�,$�6�c3��촟Z�~��
���d��ㄻ�M՛"�?�~�:�w�b"�x(�$�	������K $���7Zϴ�ynP5�.d�����9�E�0O6i<�����GB{s��cqft���:oa�+B&&��>EJ�A��9���p�,p*�0|��?�ƺ��G��04ɝ�nHG��
�ϐ�[<���Ź�I
�U�5D�k��e���!�����#0���f!P��h�U��K�xTo{����_�m���>Y��v��݉��w;U���Aw�Q����@�{@�@��V�[i��=������q�:�Y(FNM +�مq{+7��_��Q�<���-5?Pa��k�hdv����Q��k���|I��6�� ��TƟ���ؠJ����򹊩�@�L�`�������V�G��]"$�	7-lQ�{q?
ZUβm������רu=�PS�%qs5�?BA�մ$f@�Z�Bq☘4)�:)�sK�0ȝx٘�BY����"T�5#��bDe<�f���]�N� _��1�Ed��=�Τme]��ńV7�	�h�z?d_��t�}r}�~�4@�<�i�t�R7u�
�\��]�F��������P�p�a�1y�'	?���W<��ş�qb�H�~Њ+�#��tf����!�+6��8K�����5vG��L��|S���T,�f=��I|L��u��j.��U	&��5ƛĄ���K�][�L��&���p7$o\�Sc��̸��c�o�P��uy��=��4$i��>z�����^��Itv�6�}�ҿ��/ֿ����d��J�Kq�"K���������F��ݪ��$����2�{�q��~�2Q�=~s�o������ r[�ڥ]�q�X�oG���{e�XNn8M��uJ�?�tcyi�v�oO��¹�z���}��ٔ��V���i��0��i����OhE�b2�9����q<wM�d*J��"W�6L������~��AH���V��7d!S��=\]AlO�|ތ��V�-C~������v1tI�g���m�4,�I_*��DЩ��J>�<����v^�x��k;�a�`m��q�~JQ{/��YX�3�����.�d�)�w�y�m�Y�����n{;ץP/[`*�j�e�[dͬ��n߃�P�I�[��J9ل�"4^�Δ�V1a$~�y:�!tل^�+�G}O�����VBઊ1D��6�<��_�rImjα��Z�6�2���s��d����08�� ������Ao3�xv�g�{���R떩��k�H��<���Uc�*�[��G����mF���T���V��HǮ���]���X�Iۧk��,�D,�����2ӫG���x�f' �{���phRF�纎�V�����4ܣ>�����y�e�%~�h�#J�B��w��dd�$0m/����Q�:~d
|I�ꯘ-%��E(r;{�vϼʹUA�����v2�j�%�tdεrVD}�w\�P��m�O̲9��������+l��4O4����).A�O�ʨ2�d�V�����%���)��͔�@�a��W����V���т������O��J���C@���H�GF�ʰ_����X9�����/� ��,�ݲ�28�yڗ���ř�?���������DEsg��N�9M�Y�l&�VD��Cv�K.�Jl��
�Oei���gK���tS웞�I;���a����Qc��M��ҩ���厛&�
�as?�d���	Nd�N�vi�Y�0��A��J
�?\A'��������;26����;���p�tW�f
o�B&��Dɮ���](����J�-7�)�,]&o��*�Vk�o~Ov��+a �o��Q����*I���W�v+��&9xK% l�L@ �c}�E������N�6���L�a?�P���lU�dǵ�52+�΂p��s���s���f�463�,TX�d��;JA�7��:�y��S˪�eJ:�%e�xf~T�s�/�.7��!_L�b��J�1W��P��o}P����NUdd�!]��$T�����ؾ���[Cz�zd�hU��?}K��/�NB��%-���e3��dGcE<�K]բ��Xq�����
�����6_FY戮Vcx���,>eW�PWؿ���/٫�Vה~�7&ܶ��Y�����~}���v=[4љ��Qe�I����x!��%QU$zaO_ᢉN}�;��2��o�����Gb+N�ͬj�����hM*]�$|�T4��l���X5
r����
ul[!�wr��G�e3��9JqI�&/�@Ǎ��U�Pp��7�3���n��O�Oy�;A�2yb�ؙȚ��� 2��P+/
�L��j���6-����g�QR�����9l=��v o&;�.6�I.�����8��%OB5$��̸ה����s��&�D��bK��$S���ׅI�|�$9��gZ��T#�MC�]�TV;�s��L�2��&j���3�*��%+�
��{�9
�$R� e�p��6�m����,V&9I
,����A�Uw�i��3��Ǚ<�,��C��eoۼ����&����7������c[?l���;�Y���5�-�2�d�'H�z�Y8a�j�)�ЧE��4���(Y�/`p��L�/ۿ߰���|�f�̉�o�ެ���h�8n������*+��`��F
���
��k�S��̪.���O<�-�j4��틚�Bݵ�Z����������D��1�݊��ZU�Vz�)���3}ie̵����Gu�,V�g��:�5s`fE�B$4�^�7� ���<W�9

����?�X*�nAd�W4��l(Qb���Slv�\�G&����D�'�a��d>Ɋ	@���q���X"}��$�π��]#]�i�ifK��zC�jQ�j����/�}��:f�(������Ѱ���4��Fi���n�đzb�H�GN]�fu���~6^�=*�dql`m�N!���ѾS鄓��y��!jՆ��Y�tg�Ս���0�y1�H-g�da<�j�ڵK�0�}CdόH�C6
��8��e���l[�[��%�x���k�a%�7�R*�4�(VaO�x	*y�S#��Jʄ����d'��V�{��} ��%��zRcp ��K��fN~�nҏ�4yPRU#)�4��+�X�ȉ��u���� �v��e�H�i@@�ߋR)�h�a�(���,�T�� h��2��?L"g����y�)8�������� �"2�ae���?Fr0�Mg��:���@K_c�-���x���1�+���>�Y��x���a��R�<��(��>�r!I�������R�m۶i*K 1];�S�z`�A�8�#-!��3�A�I .΅�"hp4"�q��=;|�ˎ��0������~c�|�JAǂ{��+��_E�S���0��c:b�V��1SN>��|rKs%Բ�'A��ۅ��Gsa���u��$S��Q,c��(�o{ �ɺ���������.d�kR�J�&�* <�W֬]�+I�T�Y�e:�N��6Lą����49� �7�t���J;���I�6H2��x�
���l٢yG ���q�NpEf5`�ܑ���p��\ԈfYKm�93�p��Y	��[��V� �0���A�i,�<l�
��C�j�bH���D;ܘ:�h�ΔL��4�������������c�DQ��	q�r�~s�a�<��%�Mo�\آ�7r�,\��;��cTǅ�1��;'�oN��%>�N�dOl6S����8]KN�SsS]-)���i��?����SH"�#X"�Ѩ�#F놲|����4�Zo2.JW�����SU�Q�*�
(/ѿO�e���Zo����X���C������?�����,�d����N�����Brx 0���&�s�� �6lP����5XU�"bsu�	��Hb��T�qR7)QT2�pT<8��Wi�`��������Y�eX,bڡ�x�k_����.���j쏥������yC��]� �u��cB��P�z�pH^�j��?�fy�:y�O}Ɯ�,����D��G�AlݺE6�y�a�k�I;&���-n��<$���+�V��ɌVӕqN�Ľ��%*��W�xq¼�H��O~_��H�
�C���[eϋ(1�0��eX�[��+��qҭ \m�һd���i�݋�a�~l�TO��o�,U���~�µW�8V�� �}�k�����`mJ/�㔪P|�����Pc �.��'f0�0���Pc�҈��l�����0G]
���|��s���8�%?�D�
���ZY"q�h�0ox���V۲ap 0J]#y�\����Z�!�g��i�J�u+��f�������xg,1�אѡR*�Jo���3f@�W�W`:o�T���?W����]2<tD
�b��j�>��P���XW�f0P3?����f9n�9�d�n	��9X��K����s�>��7� _� H�նo�A3���yC|y����Γf貔���19|��3�ʥ���A�b��.��K.Q�
5�����Z����K�@LLw�xu�ʀQPa��ΦƤ�b;�(�3�_y�zl\�#S�� �h�'�ö׋��nh|�%	�	�7Ζl8[gB�da>�.t=hVN@ðq�/����P��-oy��p�z��䤑M�n�lT��E���n�]�xܑ/<CN[{�T�jR�c�2&=�>	¢�A��w���$g8����^��hr9�%��#��NH�qQft��.��Z��J�]��ǂ�<Os^pS}p¾]g���s���]ق��Aw�]�Y��5	#�T��_��������37](=}+e���%�sE��Di��D����*���7�Q���p�
��&�^�O�N&f�>q k�@�Ŵ  vu���0��ׅ���،�f|��ya��R�to81�
����v^0g;���1�`���K����R��
2b�ep����s}���	�~pTc@lc�Y��KSy2:,���o�CG�w\w�|��~P���Uw�-[P��S0��]m�!�/j`�����5�r�I��(@�����c���5'����QvfLD��ᩤ	�%��6��d��~>��d��Ȁe;�f�
	WW���b�D(�Ұ�;�U�����|�w�I^}�:�$n���:2��1B�';T����'� ��xF��o|C3�x���cB�L��+-���4�j3^���s�9G���.�/񼸨n�q%3љW.xիe�V���͢��Au ��2�=�VFZ=q�`�X*@O�

�y�# �����1��� �=�EB�C��&�r�3v�z�/ˮÆ�#׾��r�Ƴ�H�\�=�R�%����*�&�M7��?�>�cϑ��X�~!��Z�Ɯ���L�)�SK�|��3��ɖ�4�C����$66PR��(�hE��|*��'�#C��� ��������o���$\Q���B�%m�F�9X�|�f��gT�|vK"F}0� ���C���j�ꆁ�Z dۥUki���QË��0 j+ �m�]gc����0�#D��GG�sww�,�]jf?T.}	����&�B#��J�̐K6&����� U4uv��^`� o4�u�E)(��`QEóL	�aG�Ql�j�բ�9G]�
�ɞ���W�R(��q�v�0`s^YC>���F(�rA�"��Ss��2�R3$���F��o�'ʼ�� ���V�?��@��/��� I��]� \N�1*���֌����<E=�4�����_)Fz��PS�����N8r�5o��V����~����2��GU`�����) _���f׈㱁'�_i�L��k�E�8p>X�~�NJ4��ڌ4�m������zG@�~\r<m$���u��S�݆	�c��ƺ񼯶���C���vyp��1C�AXN��6=�e�#H�9n���`��=�Z <���F��$U���h���իW�c��_UU\x��rҼÚ3*'��4��1���m��ҩ>�^I��7�Y��̘�4OE��(�N_+�����^Q���,�*�d���:>��
⌗%S�5�A'�|4��+��B��?���`��ַ�>���W�E��:^ ,Vʬ����	3���������ň�^���o�G�Ŏ�B�2Ci��P�HB�CC�T�uȆP��#�^�3o������6"�p\g^,;`�c��g��n���m�Ш,�d�-f�p�GI�RW�}Ǖr��uf�#f�n$���<z9�!mCL.���%�񔵬BC[OOY�v��r�]�I�5�4&�=��i�3#`�
�&|V*�R5P����w�m��,�l4H���"�5l�>�� p�+b�R�����a�TI���+gd��{�n�u;Y7�0xtl�f�p�+�&�rF����l���0�lR�,�	І \�6��a	�G����+2�z-��5E�Y��=��i�z�5[^�.Eؾo�R�a)[�H,訙�r}o./s�mFiƒV$B.�J�,�l�X>�W!�����w�������a�:�I�/pF{���p��+u ߫��Zə���L��u�8�]��.�i{Eثvb�]�3��ZT�;n��av��f�d�t�޽gwa&r��s��!60c����KVb��	t>X�}��j��1z�3�ZSt9a�8�l0�x���L��k�&kVwK�ё�ډF���U��w�j v��\rɅv��h]B��a��H&���W�z�&9p�jƴ!l^��ƀk�*X@�c�Ft�}Y-dpI�� �|���U�7���M]/�����`a%�&��z`K�P�.��L��8�N^!6�0c�ho���%/�̉�����C�>�3o�G6k3P���8#��f�t	ܴ��Q��.�@����/�J�;�S�>h�d�Ri�hJV7��Oh�=/Ԥ�1�kʂ0��D��U�ȴk�I.��,6���!���c0�oɀǲk�a�f|�1y(�+A\��K�Ы9�%�&Ԣ�H8dU�v?�3�~��o���b#F(1�0���hP&�5p�2���`/�ʳ�C�'T�����̰�l�A��۱=NB�"�v��.v��e���
ɰb�e8�<�����m	�m�C�d�� t�p��<%�����;��N?��׿��e$62�����3�f�.�8�!��;����Zal��e��r���xE�D����9�����$���1|ė={�����ʿ��0@\It�KVʅ��L6l�,�jA��T��	�1�`E�m�ZWo+�(`��#�ZU�(�*#�@����/�O�Se� k����A= �
B�0�wbڝ�{L�>�1��X�Cg����Q丵�/�Ӥ=H���i7|�Sdͩ����v�B������22[l�9TS4
|�q��)�/lU�*h�x@sV����W=0ddT�R�����k*g7;zNϡ�2�z���{�,)���dd�%ʽ[oאK�)�z�Itù��r��a�a�xH8f:8jخY����1g�UW��zVv�8"Q �.Þ_H��bdT��.��	CM� � 緼�M�w�K1��f`�ƍ��g�����4M.��{�,@*D�­1��< )	&���`b���1���]
ޭ�֧%S�@�q���5�46<�����Q�W���iz>���'b�`���@��D�!��@��Q n���xȀ��׽N�?�|M������w�yg�˂�Y>L>�l_G�(P��Ǝ�&~�	{w�'G[��I%Yg����r��bѩH���c#����#��`��}��zV��L`G�B�a��ˠ��/�\1*	�{�W0䫮z�zI ����؏!�XM�}�ٺ��k�y��3]Ѩ"a� �
j�B�rg$�Ŗ�����W���a&�)Kr��ae�o��W4�-"�1h0�0���m�f��@( �3�T���x���q,Ap|���~�#�aψ£��A6��j�v������M1�tH��}�谖zA� ��A��9 ~�J��\��j"����� "߬$R,��f�r�[����%W	Md ��{����1z��3�Q<A���J� �
 @�E�[F�# �XK��X���Z�� j�0#Ѓ j�'Ӌ�4�[�*�xܡ��ry��u�}����I�q�K��0U�/]>(��|��iш�1��64*��P�c{�xA�ш�1�ne���́m�5�|���Z��m�{��#���Tmd\JT'C��K_#KJ����J�����{�O?�9��iL�	�{G�KS�	M���e=����͐�-j�� h�#�[jcCK�s�Ӵ�fm>�I�'���'O�'*K0h؞zz���茡� ��ؙiob p� `#	��h̳�d��c�j,�+o�\R0��EѬ�x��	 CK�(A&qs7�x����4�%t/�@4
@I��x��2�)l6����l��m�+N���ַ�_��_u6�;�� �i����m<���MA�v�5]��W֟�/���R�nؿ����zc�lT���@��K./S�ll1jۙղ?"�#��ϕ��/5�-�Zݗ�%�dhDd�Hu����%Mx�[(��N�8�˞k@ژl�bF�Q��>�W��W�{���El!#F�3�[L� !�*$�O`â������r�2%������)���Z��n����Q�)4 �?�p�P5п��@���ҵ��I�[�:�K�3-S�Q���I�c��M�����5������w�*�x�2��WF��(��1;ʄ
��
"�\�B*�]�t9R�*pT<�R��0��g��R.��z�e��f�4��Be<	�e��Z��|�{���!���R�� G��2P��f5�[n�E-��#�T����nE"��(��W�?2d�A[S��xއD�Rr���& L�\�ׅՑمpcL���7�$P%@����K�.�m�&�=C������N�n�mG�	������n����\�����~�=I�;�&Œ+a�O?�t;izG���\���}�q��D����O��/ɑ��a���/�B)$KZ����a��1�RK���$�$\d��![�1o�!h� �Pi[X/��+j�t�������F���4@8����Փ��F��t�F��(�=�ܣ���p�`��t�t�̺q���g�Zb�b�v���
�\��������O�o�2y�������T^Օr���Q��� ���AF8�2�`¹�R��x��Ы:�P��ȑ1�η(O?�O�9o��
��QU�Y�J	p��G�3)����%I��	!���{�fDw�$�D�	�� -A�o&i��JX�]԰-s���m��(��t�����#L����F�����Ibv�#��IC'�r&�a�N�v @B�wG�@;����'& 3���3�����y[���;�1�Z=���4T���!����3��G���p��cN+�%�s���(��
�� %@HT߈Q�H��=���o�A�8��B�*w�X-�4��G�=�EŜ[�h����e&ۡ'�"@�`l7��x��A�q��-�o��D���t��'�5�ˊ��VR�l$	��P�	�	�V;C~z��4�����!�M'^����%S^��G�=�xiE�$e+�:Z�\���hM��ukd��^��	�F2+k�'4:��xE�"���\G��	-�M����)yAM���a)���c>{�OFd����_��F1��;�D��h�U�H�^I��m�I��u,��b�h<���`��,��[ u�+�x;���ΤF�i��m~�#�:,ms7�RLg���Sh=���Ͳ�6�O�lp���.�ț��Z9}�Js�5e�����ۼVPȓF��rѺt,����%cY�r���(w�����0���+H���t����a�Q�
ؖV�7������*�e���k8���m�4 ��m����i'������
Ϳy�������W_$�>_F���oH�kn�%%Y�AA]��¹��2]7K��g����Uv|�����V�%�Ε�����=�<%�m0+��`<�KO�Ig�
�)h�iE�:I�l�j�6���,�-��`ʻmwޅ`��9����Y���r�\w�I{���kd`�82:�G�{��F@Å�HZ��UU��Ē�ͽ$ryy�L�B��s�(��q�h.n��W�s��^s� w�X���a�}�[8����
3�b!d*�k�UO�U��pڗ�H@p�}@a���YҨ��&���hp4/tɮ���ޗ�S��}���+�'}��_;��b�X�#inkʼs���*���o�`�R���3$�>�TʮV$�`��nCnP��W�zz*j�����X,5UIƴ��I:n���$��L��|�$l��C���eɁ&U�hؤ/?���Q� ��G�J��%w��7f����J϶ *�\r9f��T��������/_�Ï"��z�R����.����H�>f��"�_xN0G�1\ՌN�Jq>e:㺵Js���)��Ubs�l!@��jvA>Ɔ#���5�����ȣ�J����+���74K�����D',	�p'�c8�8'¹��2�N؝��Xj���Q��P��[��CU9rpL#��9u�iV�������Q-�nV��Ɛ�m ��u[U���e��j'��Pf���L8.��G=��[�k�B��;�=�Tn.s]6W�G��U���=*cպ��`44ܐr�Wg�(4������)��șq./_It��JQr�a�%�u�ZS��4�;�P� v����n� �u;�-��خ��v�9[��h�ߵ��>w�I��LY�PD��$�,l$��+4��&J�-�I��pa���Q&L�l�윞�R��J����2:��˨��<�s2u��C��X�A����eI��3�_�¥c�Xv��oZ�dfq��S��d�K�z	Cfs.����
^B�ό���O�r14���{��J�Ud����s�շ��a�F�s&c�d)C�u�L�Ê��b�[&�aUb k�� ˀ.������z킟�1�EG�d��$���a��1{zz�Z}̀n =�.xhHZϭ�՜�ņFBR�(~G�
�Ff8�^D
��l��j�T;п��!8/R�m۶��}�X͆-� �cr�%�ȩ+��/c�vH
^Yv??,���#AL�k'�aU�\���[�	���<(x���m���_s����(�����JWπ����@���$w�nB����Gi����d���$��l Z�s3�Ta�c��8����-xEl���W���6�+�0�u��o1��3a���&��PNA�4\���(�(�2�#�rc�b�ID�����d(�<�c,�^���L��kց�I}���=��v�{v��Y�j�,]f�����e���X�W�è���!륯p���2�U\�9Qn�w͊�e��+e��k��2#��,�{�"8�l� �w<I�kV���s�	��I�ƒ��E6��DJ\֤c}8V� p�եy�H��w(���cH��c��"��� =/����$?�b'���E;˄����:�:�r����~
h�,�����9���N�c�[�7��;��s�g����Td3_;��L�3����s;>,6 ��m��dQ1�����|�;?�姊\y�y�Uꑣ���<ui�m�M������Aƽ%�s��\���
�7 ����i��C>b��3r�+6��ҵZ�hp`�2������Wj��昧j�Ł��^�n���oЂ�x������T�A�3���F�!���r�RG^x���e�&� �ׯ_/7n�ԙO<��w�}
�L��4���0���.��eH?WR����ޛ[z����Y�K�}E��,�UHB�Y�&���ej��$q2���d<N��$�q9�	�+�8,�)��n��lV�f�EK��u���Ϲ����{���,��=}�{��Y����w�+��x1�����ԧ>�0av:���ݽ�,(=̗]��{�2�=I�u�<��:9��9dÂ2�d�����`�u	|F��]�I������ҭ�}N�շ�b�W�SZ �����56PE-�k<L�n?ŭ����LZ<:H�ƽ����|��7��[���q3����t�g���n:vl13�L�23^�2��U�y[�l��:�x�С��]Ď
̴w����Jԃ	�b��|!��`1��Lވ=���ݟ��g�b�A���1�y��:��p�ȌwRQC�; ���W_�����%5��vJ�U/� Tt `L�|�/{���������Ed�2Z�������M8�ߙ�]q�tF�s�F��4�ޕn�w)���>�^�ꗦ=yw�͢�5҄�6ƻ^1F��~������=>6���o���{aW�0:rd9}�K��y4��}n:�A��Uu���@�Y�0�5��0w�za ���//�-�+l5�ھ��o-Y}-��|�W8R8C\��XU�n8U�w�W b�
��`Zވ��q��B�TuG��d�3���b�W\�b�B'���Zn�����+��F��1�bԀ#�]�a�9�
�dԏ�D��3ϝ�nF�#��i���Ӓ��V�6G����#���=�Kg��V���r5t�u�J��ԛۮ���%������u�f6"��jf��↶��F����%(������{~nO"���)������!zW�L)���^��������Zv�.Y�^ı�_�����fS�hZ]j�=צ
�R��O}j�'~_�3��ߜ&�\cm�
 .���.�����P`[r^ r��{��ǘ/�݉�s�}hV�P���k�413:">�q��Lci�%[�	O�y`�=x`!�����w�tɥ�(;�m?��T�^�P]5��_i���"��On���V���[�A:ppoY(`��$���bj�T�r����`�a,�{�����׿>�����9sPi~��/�(��z`p@�<N�9F�� �O�g �#<ª��ک�� �:a�Ӛ,hְ�o~�bE���������Y ZU�_��إxO)w/��ӹ7�x�D�s�e��7��嚟��g� V'lֵ뷊� ��j��28�<7;H��ޖ�>��~�^�'P?�:�i�5̬??�p!��$�ο͢S�-K.��1���[�Sth\��}����y4@F?m��ڧz��rQ���vjYԪԹ�"vI��F��4�8��L7-�׿���;��a������j���4�5J����Mb h�8�=I�UJ�ˆ��R�N�Yi��S�?%D���h3��*N~��wx_�)p��7��#��qb�y�0����T�h'l9 �w} :���x4�-�-�8�-��~����78DQ�?�y�+�Cf�!�}�����ɶ�K��H���_������M/y�3�����_�UE��'C�U#�;���m.ޗ^"�lKL��;n�N�h���X�Dd�n������T��g����\��Y?�T5~B��������矕�ߟ��|� EY�̆���I>p�#�-O�w���~����{�-	�N9C�DL?ap�ȹ�Pe�u T�j'�JǞ]�I |�q�� VQ��j�Ӣ��6[#
����J�{��Ep����=g � K�U��P������b{�7�]��r]�Q�����¹0���������ƸX�^�i*��p9��k^�Ͻ7ʹ3+~�<8{R#��=��H�J"�VI�<U���$b��[d��h=K44r���T�	&��]<z�ȸ������v�"������n�yN6Rg���؎��/��@3-.U���>Et�ra����*��!w�|�+�}�J	 }��^W�v�3k�H���Z*�b<� ��wU1�.�<&�%�h���[ �ƹ  �����������[�R���� ޣ> ���}���RA���*2�XE���y���<�$��KGsM ��y��P:��a7b `ٺ�hԏ/zD�VTX�,��XZ^z ���I���X������{�M�Z�8o ���/"ب(&��bM��m�yy.&o6'�);�`����[�IVϹ�eO�ux�=�N�� &��4���L����a/}�ۇ
�Y\^���@"�e�f�\�>V�N��M|u-Q���i<#����+��+��ha� 3��,�b�DW�6d�u�yX�ϫ�W4*y�5br0>7�x%�Vq���ye�~{�l��t�ܗ!|�H�´���d\��bu=�N����C��DM!0�.���v$�Gv籜���ă����u_��O�E:�A��]�b�L>W�@{�(r$��%Q� %jy��K�V��ʸ����E]�j�0T5�*��=M5����I����C��Oг�Qi��Y�}���p��jYXN]j�5g�����@��}��<�������ԧ��g��IOf���	�B��B� ��x	s� >��a����// Ѹ��_��_M��dòZ�$K�i���un�cP��u�߰^ū`��5��'-�@�a#:%G�ca����]E}���g�C���9�������i����.�@�f�
��`��ǃ�q�tǝG������ئR@+���#�	��E��䩨� ����ϝ%��z������"Fa�EdZ���u�ұa��i�}��Q��jUE�#n�ކ��M���`���@:� �Ġ����N_���Ro8�v��W���Z�J��5�m٩�8!�vQ?j8CB�s��$aF�I81V!��=���ʈ�bU�-%�9SU��t�[2a���1��;�t�X��JS��aEݬ��q���*������s?�sE����u����I7L��9 !�z���q�U�5h��ǎ.�ߙ�T(�D,/̏4d�͉��N5U'�!�
�'篛�����T9�хq� 6�kâ�@A����n��i���zl5W�ˣ�l:�o���}�53�f��i��+u{��U%s0 ���s}����%����__t�	� ^��/�B���K_��d=�*+s�|1߃8��*=u2�zL�w����T	�����fba~��0&x��߰LK ���/ܴ"1/:��A;Oe9a�Oy�Sʵ�h�r8\�{BC�=G����c�V���y9;w_a���ZNS��}[IeY�n35ơ��;�!a߸Kc������x={_3<�Z���?��	�vr!��>��p;�&s��0�ۿ�_��0��]��G{i���+���t�y&\������'�u-�p�*6a�Q?|�_,ċ(]���[��������19�	Ŕ4M,溚V�^���o�h͆���j��R�#3wX����������V�\X�5�!��%�_��&��:��"2��`��À�d�X75��XIaȷ�r�:�4�2p:�n�����b��G�s�:����k�]�9������/�M:t?.xc_�̊[�,�dq�2�<=����L�i����y��18�tD#��_c��Q� QU$kv����Ltth�5.zi�&��w��=�L��6S���XF�@���a�xhu���UWѥ��t���$}������w6��ką��&k"\7�֫�G����R[�w�1|ٙ��xo��g��y��c
� �|��a<�V~W��.~���RZ��I׿�����D������kj_:t�r���嵚�d!���R&;�ɜ0��}��������da�>D�џ����xЪ���b�c."	j�S"�?d̮9��\�:΃m��a��i��= �k�
h?��9�Fg�ܕO(:��sh����u��Iv��`���>|���$�G'� �)�n�p��x��_]������c_����{
�}֞�g�{ݖ��]�Ϧ�G�������q�S&:��V)-]�p|��8X�N& �7T��G����*0���,��~LT�i��B�A}����P�'i�L�{=>TU�QF�`��p�İ�hP@���gU/���	N����9�*MP�|���Q�V/��-���;�s��ϣ���B6E���e���ܳ)5����s�-H��<����@#�qv�H��;3Y�휛n�클w��|?���᠚�s��
��b_��hyȚ}e�-9�����8��:"��+[UltWaɟ����٫S�
��0r�1���c��K�诺�:b0(;(*�Fw5��3������Lam_��m���{'l��N+�M�/
 �VIgG�'�k��==' ��Qrq���:�I�Ȼ���=�%�N/}�uU&���|�_|�+�
�K�V�\���aqY��|���	�eE���=�š�Ɂ|�^���|�P�[6����~ٲ#:c�����S�]�)�9�ދL32Q�aLQ�u����q�J��#�T�yd�V_�Y�z�D�d?:�K.<w��7,A<J~e�5ת��kՃ�di� ��IdA?�d�3Οh�	� �5�'��1�W��x�H��習���;��u^c��kj!�3c��0����qǹޜ�(j4�o<�)
xUn.���д��է}�[[,%%�$��F����cc�N��a\H��^͋��΢��b�˼�E�/��n�_��0��.�@B�I�p.�n�ݜs�M硎` `����?��q�9�~��	 ��3�w��?������w|/���ki�����x�̍˸���p�*�{@�G�υ(D?�@�L��������6�}d�ѵOp��h��Ah�4Y�b~+7(��5Cb���	�Q�$0{?.n��D�n����5Q̶��'?���JUo�%���M�׍ȹ%<�����_�ӯ.��q������� nbq#s�� 7A��im�0[4r���Gy�U�����O}6����p��x�cӹ�<�����d����_�&m>_�SЇ��<�����@U'@�o�1@���ߙ�V���{^�_ԅ`��h�h�9U�bK��r��
��Ro�Q����93]����	(?���"�
]���O �u��7�u�v�s�5��l&9�'���an�=�9E���6l�Gü Wf�L�t�Э�ܜ^��Wd����n��(�bW-3qq���l4� �lP�0h2w�v�;��0�3گ�GH�=/}���t#�n8NP�;>cK�^9�qa�Ff�y��
�W��2�"G�vL;% �G��q�,�MH��8u�)����5"��ܜ<FՖ��(mE�瀯h0�*/��>c�37P����p^���OfU$l���Yn�;����,U�;��̀��S��?���L���� �H�3{��oHވ̀��Zq�g&ܠI"�wr6��C�;�L i.�p��Z�7S�!�W�}�1�Ҝ(�ɑFh4�K�Q���Ǆ�����ԙ�&ʰ�ȳ�FH�������9(�n4��X����R����\�1H�΄��Q���
 �~���0,7B��$N�i�w�f�4�.��QZY��zG��G�^���Q	Ψ�q%jn���ˮ����7�'�('��G?g�&��)�9�A
pH �}��|0�H�'Rt��.:���rl�L6&㤟�`6���`4�����S}�s�0>��0|��F7�� �|�����I�B��'HMH��ؐd�qSQ�%{�) C@���Z.���/�'j07�>ᚑ�sN�ec^k�+�����=��}�	r��n��e%�Fȋg�3���X���^��X��T��d���֓m�R�;@������R�mi~�=Q!��.�t����VW�\�j7��h�q#a���H+lB?#�b��ߌɾ�O$k )�1`��r3�|�K�.k�����i���=��	�pY��qb��Z$7��}�U?_��xy��ޛӏ��C'`���V^���O��ѿ��22u�V\U��.�-�.5���#�o��]�1?��47ߩvw\�y@�����]|K��Z�Zd�47��X#��%�3��cq�|8�`��=��b���5�y=@�	���sr=�'��1n&61�}��pO^܇@��`� ��K��T�6�,����*�(F��l�8�RB,�8��3D��碿8 ���>�*��d!r� Td��C�ٍ����FgF=;cʼ�xv��k�q�A�����Z��@|]��+7����^釾aL7�i����y���u�hlr|��V\c�H�ֵh�%�0������-_�tZ^9��W�TV�Ro��O%-�Š2�>��������L�N���$b�c�}�ܠ����\��܏���S棛�7��������4���Ä�P{ǖ]v,B��8=3��;@�A1؉�Z���� 8<��� L�2��������X��L�]�RGk�ĐBrZL�ѱt���k_���o?U<�٬�y�\|���xK����c��+�s��Y 0A<;;����d�y�(3��Ȩ��::`�o�0��bԡ�W'Ɏ�(e�dt�������E��Z�z ��4��� � '9�x�\�  	�`��Y����8��XO�7��H�ȸ7�ɴ� ��/�ʋq�1�[�+�2^�J�^\����Fk�Uf)���z�2q>4�,�v���M�f�,}�Z�J����l&|��������D���jc�(���u���^���7�Iǎ�*n��3.4Y�_cCl��h�`�C�����9��l|�w���*PؠKQ�<2n�ĺ��2/�|�Ӏ���uPI4OGe|�h\�����a��Cgk}&�{x ��i@Y���q~ݓ\�.VZd/��5�e�F �<��n�X�巼8]x������4���.�;+7"sX��D#���a��g�0� ��A �=@�Ŀyo Qt�t�@�
:��d<����u�q�0q����@�_���7@������)++��α�ȸ��m��c��
��: 'ǨnBtw�	�	�@̧Ap]�	аy���>�=�T��{�ч,n���o,Z��A
r�`�m�9�
�G�c��&2�ڜ�{��$����w6#E�`4P�M��J-�M���dW��#1���m��7��1F7S	W��O�Of��
4�:�t��OM���_������ݗ�^N�),���3�ɿM�յD8�$9Gy�����$��x�zt���s�����%��8�W�	c�ԤD�9"f�~��eW9�v���'��ڤ1�&�L��Jv��]}��.R��04���N� �N�\����H��ufK3��dYJGg �<#�kp0�1u�<��[�d��hX1����So̱.>����j� ñ���KF��FR-� � E�n:>���cf�WU-<L1\�~���Y ���L AF
�D77�Q��T8��D��F]8��Y@�X� �̒��&�Qm{���g�"�2H��	�P��Fù ^���D#z谈�
��G>�w>3/�~���s��K編 G�����������@�7� :�W��Fǎg	e����=��I��{Rz�eOI��q8�%(� ���u3��z�5{�@jڏ<���{�n*V��Q�F��-~�M�괂���r�Y_E�����;���71Z���X��7ͤ�c�<yVґ{o/,xi�P�`wםKiϮ����V��-�T|�["�.�BTsL��04&��� ��,� Xu���H��Tt�R'U^[�'���ٟq�k��ا �WG���ʱ��\�c`|����s��Z�Z�#(��k��Gi�DyY$ �U34[=�Ϡ�@����ʽ�QﮇC]�eC%�􍢪9@3�2 $�����k���`7�=)��F�8+��-�:D7P6DI���0�w��\^s3�3qٗ�{9}�����9���RI����!=���46SoP�0X�������h�٪m���X����<Y�:U���	��E��J���^w�W���xF7��4�I􈀙�K���.>�.��|��t�m��UG�u��ؗ~x0FB5*�Y�k�=K]Ɩ����+�5	\,,,�	���{f� \FE7����䥩/s#�ݱ��q�����
U�?�������q������ת\x&�	��S]��e�����P�%����iaG��Ёj(� #�� r#]Ԝ���mi����2���ߨO���@�uݬ K%#��|����W\1�ce�@�õ5������_�}���;679U{���k�ԯ3sԞ��J?����P�;�+���l6ͥ��=�Oyj:�����-�O�Ae������Q�3��~��\��8Y�\��hC�<R���g#p>m�9��6��Uҝֺ]*�������؅, ;�X��3Gv��r�{���ߕ��⢴�'k���8�5>n̂U��kTV��+�0W�A+J+*��M[ɱ,,U�|����vk���;�"��C���T�D��!@ �y�� 2T��H�� J�h��J0�����Q�j?*N�o��c`��b� �1�9�}��9@��M��{�e�</��Xm����,un���x��Ϸ�0��o�v�zэ���=R��� ��g>c��yO�rO܃���+����mie�xu3��ՙKwޅ��0�u�iiq%s�,��D��_M_��;���O��*�Oou9u�k�ݴUD����<��u+6IQ}�D�9n�_�P����V�Ś_��q*t�悎�Q[�f��j�	�R�ޏ��Z9���n�ñ��ư��2���x���ΕdR2��;�LD����H���}I��E	u��'lN ���Ɇ]��O5@�0Ѓ{U���q�����p��waEi)�J�� ��|n�7i�.�2{p֪���N���e���Pk �|&+���>��g}J�����oA�<ԧs�z�"�s���_�{g1���G~ �㬑Q��:�is�TZYi�@�k2��H��k�lg>=p�p�x�ymeIs�f����q뭩H�7S�P��dY��{^/�;&1�cں;�6<�>�j���CٱQ�w�����hQt�܈��)z��]���w�?�>��v���ۊM���͋t�'}����ˮT��UڞQ�r��\@,���F��K�]��_�{ݗ�C������{�u��g��M��GР}m#�	���c�e�@�H��]XV� �Ȟ�q�Y�C�X]4��n�V���F���7���]m6*���ٜ 4@��ͣ
�ee��*[�?���+vC�9�q�T��=��<�c�}Y�����97� �q����g��8�\�f��'�u��%B�7���AZ�k璟ɛ,��a�V&��iqeX<%�>;o��"�s
��5Ɖ��/nt�s�"^�}�@=��u����I�N��Vmk�Q�7�r6��Q_Y7Z�p�e�N��q���Rv\�?J�P��ꫯH�w5��0ͤo�ݽ����+--c��)���l1QRe�{���X,�7%I&&��hp�K�j�c�O �jl
?�:���M�P�F+�6Lӭ�H"��d�|�ƌV�D�@8q,L̠��	ȹ��Y�d���� 2���Or��{�J�O�HI��
2Ґ��q�:�ܜCC����;�99��bf�������a����>�zƠ�յN��^.1/�sϡ��q/2f����y��o����d2��F�w͑�}%�⫟�^�����\� ����F8+�uj��ހM4K���q�8#Q�g��W���؅A��&���}��(���	��)u� <�'Yv�F{,���+���޴U֣�L�"���Ț�nRu?��8��1�W]�_WV�r4O�t�y{Sp$�u���{:s�U�fv��"Q����Y�k��i��gq#�i��j
<7� zpO�v}!c�W�u��b�w@s��Ⓟ�j&Q�xt��h����LQ>NJ~g�f܀��70<�w��ƨ�t��i�y(�4�Ѧ��c���{NXolO�1X$����iج�5��|��i�IT�9��3�a�ul�;��^ �^ݸ.���q�D��g��v �����!Qo���XIg�1����J����=���'�o#ϫQZ<�(�`��crS��~�n�]�~oJy��<�u��@c�*?U��,�����.�{��%Ap�E}��w�G3�^�1 �{����w;��0���F���#��ZlG���zb�]`u�v���2>]��M�ڠ����{��(�w�Bz��.K�����Ky?�J�'��+k F���*߽U
Q@@0S��ϲ�Q<e�I-�ɈQ�b�f�p���Km����n@5`�-�u"�J}��o�i�z�&���N�E°�wu�����7cqu2�9N��bۮ�9��4:�ˢ�k}�5��G�l�C�ޓ��M�����Q�yZ��G��j*��T���&��������:P�p�W�e��m�=��m'&x���.^Y��6�����:��e n5�A�hI=�və��	�Չg&"y�v��w�F~;�,��h�(6hx�^W?΍�]Ռ�O�G�VW�Lo��^�~��^��ҽk�;R��0��󰪶<����/���K.�l4�ϚU�{dN���k����0����������2�4���߭�[\ [o���������A���e�ݴ�nv���u�'�L��5�	�H���l��¥�L#��|�ӟO��ޑ��I���/K�?[ x~>��X&@�����	�/�wd���h<��� �$��c����mc�e/��ؤ�9�!"��6a�m�j��G��(�ɮG���&vH��d���F����n����=��\tx2>E�1�ц�H��L��ٕ�{)}�c�~��ǧ'�����xHL���y. b���,�Z*�4����]��x��x�C쿸����"����xYr<W��~Rډ��F`u� 6��nv���Zu�����F`_�~��6z��4��U�l���0?��>����wI��L�=�?;�R�#HPe%]7Қ7Ud���X���J�UPۊFN�EI3�����|����͙m��{)�C;:�̄��l��`[c ��y��C?5�;{�7 �X�aS�?�u�և�
02߭�u=My�0a/�N���O1�x�:`AM��s�Y��W�����7�M�K�4�!�CO?Uي�ͱKZ0Ѝ6WG��U��F�G���
S毕�}���$�ƈ��KM}q���!=���=��6E��g������`i[�ش{8Q�?۩0�킿�4ͮm#��4��ζaq�Dm7$��Q��������3/�n�B'Kγ��[J=Ԙ���iϢ���\�+�*��Y�u�F��f�+mp����_�fTc��*��k�������;�AC�`X�,�kT)�V�Ki�W�^v٣J�E:�/���N�E��� UQ�&G1�.j�26_�-:����Ź0��c��q�������/3%z����G������´ɜ?����Y�ze�h�Imb�
�e�5XV�R��s�S�z��'��rpC�Z����^@W���&�h��3��a\��Qo�O�O�}n����|�����j����`l#��Fg;s�e�o�JDe��(DXE��BԯJ���8�1C�����׾�����>������+��h�ǥi��P�{R�^y啅0�1u�\��� 1 O�KL�Ͷ�)��v�QF�E��2��	a#�ݳ7=�Q�MO�3&��`������N��YB�2�X�Ɇ�\w׏�����p�&U6�bt E�?��?.�jb��Xbm��ĿF�'$�����^���s�={h�~�2̥����ƨh�[�[���L9W���`�L��4�Q|�( ��	}<�~�
���a�s�2���I�Eo�6���7hlv���Է��&��9��t�����O���uY**J2�eN���ۓ^�/H_���gr��slD�Ƽ�g;%0jee)���KC�;���\M!��iQ�F<��,�ɍsL�)��X$h� `�qx�@H��v}qM�#�]?�9�)XCRx�m�JH�`?�ߝa�@�/���xEz�S���@y���9���� X-���z�K^���O�tRa"zV��Dڋ����u�1���Ό���>s��6�K_��t�����yr,��ե�UP�F�P��p\�5�b��DSfu�F����/����
���e�B�-�4�<�����RLS�._�z����'Y'|*m+�jlu={�|#�矦���s3�]7����a�Zy�o�
O)~���	 �ٵ��qՕ�w~���S��t�E�j�H���
��t�+(e�x�i�z^�a��3�� � f�j�pǊ�G`��W_]��
�`m��|J����{)X��1�馛
��}�Cw�v<bn4LFX�O�9�I���?���%q�s#hS`f{� D ��l=���� =P9�ܮ����{�yt ��}(}���ۍ���"U\�z[o�\�B+U���׾"���t����y�V˥�܈���A���H��	Z�6
;��U-T��GU�F#�9$��琨_/�b&�k`�zf8���g|��i-�F��'�m�з���TJh�����ot��x7A�I����rNKKi����[�>��\� �c��ֆ�N&����Go־m�b�#�Sy��J�:�=�;_gO:Vr��t��/J^zA����b�[]=���K3}���� $����Ӌ_��w�[5@H{�;�1I�dȼM&R3�������;L�B���"zd���/6�I����a¨#���w�V������Q��С��y9D=�D���H90����t�;m I����e/+�!₺S���O˥���;jW:���F���oݖ�;wEs9�J��]�����g�9i���q��x��/c��z��������\��j��J`�d�%�ƅVw@����~ְQ��,t��ͲNG;ϣD�{��xZT��bܘ�<Z������77b�"@G�����M����F�q�|��p7������~��<W���=i���]EW<U��� mU������ �?��?+��@L�Ԙ�Ԡ$��T �%8
�dyf ؠ���գ��z��������Q�vm��M��N�Ǔd�ߪr��t����
Ӣ�0�J���������≘��c�w$���~��������=�yew2��:��ӛ�[Â��i3��a7����O~$?ǝ%yLw8 Bno:t7eY�dqk0f�c�`������B/��Xj��b���gdr�䜗�nu�1Z��_f ����l+]������~�3ݝ�h�L��T<�@�b���h���+螥Ǐ�o:��^O�Y�:k�N�
M+�d ޕ�����#�#7|*�������ƹ��O�:�y�i8GC��6�A�^%g�)"�+�>��t�7��X<;����s^I� /�����D�Dc��zt����<��#���O~r���k�{O�O:�7;��Ǐ-�7LG`y��7h�.ߣ��0�$�7�	�����s��a� UX3����ԸP�b��Dy@x�A׻2�=^,��A��[�,�lwW2J�;��z�H}���Dp��P`����cSP����CYYd\����v�m3C�N<{=�JF�/:���M4_O:�]��Cg�9�c��=��!�y����������yMt2���Ez�kϧ#�g"p��^�x����Sk�R����Өt��3aUeJܣ{Я�گ��O�_�ksx󖷼� ����rN}�G�R���g�:��F���H�@`�C�Q�BBQÊ5����L8��Q<�IfЏ8�s���&�Ao�>���6���` ��P(>��3���ท���e��X:�����{�{Kgt�����N���
�u�U&%9�3C�Q�O�!��!ї�ۣ[3�g�|Ƥ=��~q��|�I�j\b����g����1��� ���!?
��V����P��7^s'�7b�H���S������77�9,Xi�;+�u�Y��$N�y]G���:uuDQ���Y:�f�^�ղ4��n����i���k���-@�_���&x�j'�cLpϽ��o,j�c��g?��x~>ӥR�˹�_�
�f�i���4�D۔BL���&�W��6�U`o��`�F�?Z�,�,����������l�UԈ�~3���b����`h��\Oy�Sҫ^��I'�[���N��z���]��a�:"N���]>�Z��,n�K/���ӘOݕ=yw�?�g��#�
�� <J�zz��|��؜@$]��ͤ#�� �A�z�gN����t��$�}:��MR	.����3]'Y3,~2���5ZCD��l�w�D��Ѩ|�����M�fb�����Yo�Uo+uB�Ľu����8s�T��hB��L������g_���\,7�T��1�s� \E��<��5�����t�5�U ����T��?Xm�g׌^��4�=&��:JVR�n|f�cQ\pW��Q�qj	�OHQn�^1�IRv�V��Wr�iD���b�[��s�P�3hQ�Q �'bɯ�ꯦ����(:|����g�z���4�M��bzы�Lg�����-�fs>�����?�'�:��j��W���/� �Q�$�9�>���V#�d'Ϧ��	�,�v\h�?��Û�u�T�
�N��9��֯����1���T�*Rm��Ҁ C�a����H�G������P��������4��/`��be�8���h�jN��ʀ`����tn^Co���^��g��YI�n�v�����l����h��Kq��\�'�nhu�6���/#���3D�����e���7}�zrܢ�>������Q���4�
�muO�7�n�5���kV7�5��wח{l5��x�~Y�zN�ĺsˢ-?��w���\LX6L�-�V��!�b[£R%�9���ܩ��E�Jn�NZZλgcWIFR"{FvY;m���m����lOQQߡ��1�}�p�~����QT���
F�i���ТԶ]��@�o:����o@�o��
�3E�����ck &��1��s��� l�k���y�?�Ò
��ꗴ���R^G)�;�.�i��N^_�y"W�(�����̩0�q�Z��(<Pi�ˢ+�U]1�`8��e�GOu��F�K����@�3:H�� {su��5[�Q���7^̣�I�JG�@FQY@�n$��Id�E�b8���Aa��/�忤�����x���S�{&y�@�p�}?梒�w��]��G�N����R��Z,�s�3%�)Y�ƽQ�xF̬yKl�Ec@l��R��4&N�i��?��(��F ���F��,+&������i�#��?kL[7)�)���[�g�f-���5%	2$��9��"o�����N�� ;�y]3���X�Ъ�Gp�B4�q[��sh��(#&��
 f�*"r�~i43�����8�7�?��R1p3�G�/�/��/n�b���/K�ܝJ5���KH�s���&8a��qݲ����o-�qG�x/j�4��{��__6�?��?�����T��E�UF����Q�i~��I
c����j;�;ɶ�N��7��(�����e��1��y[/*���w��99�w�R6|f�Z	�X�%��������b7gpaLl|S p;_fASE�:f�i��n��_�n�t����%O&&��4d�..h�qhGs��;�����@�Im��;����X0GНi0�`L޽��آH����4 ���z���UND'�[V7o�7~�� s���Q���4bT�_nhQ�S/���@$g=p�qtKs���G�ܕj��J$�)�����.[\<�n��O���7~/����ї]����/���5���R�s��� �e�;�=�)��ozӛ���jbw�"}�Ā4ab*�[G�n-� �Smj$�����)u���	�����/Y�mt����,���=�:���ݭ���CE�a8L���U��������d춵�����L���|�L����7_K��c�׿4�y�A:T�s�@����}I<2S�Χ��f�+Y�e�yY�GЍ%�l���nH��F]�|i,D3ũ��1(�D[�}Ǘ�C_ɜ��1Y
I7Js@ˤ�}�g� ��Cp�XT�1�Y�}1�Y�OՄ*9ƈ�8/�G?�u׵���GԵI�3���CZ�d"���f5}�7�C���y��M�3Ӡ�7�h&1�RH����Z��d������Dʰ"9}������whх�y	Vq<R�D�9+fG��͚��`�5�8�n���΃0MŽ�ą���yl��{�7?H5QxX�G��N.2` �cd,�6>�*���]�c���g��GL$�	��\�>TvI]�bL��ހR~7K���G��_ �LY��~j���=UG�\�1~h�QO�99�������E ��u׶�g����bFOU�=����dT�O�G�����kxV}���KSt�~������y�K�[�$bb�� �R�����ѕ������
*B4���'Ԋg�Lj6f��Z���������轻:�\�2��ۈ����^��i�Ա�y�$ B����}��.}�Z�_�7X1�d�a���9�:s3f���/Y���4c^���q����Ou[;��F�q
���L���z��x�v����M�f��e�WUh�-�����>P���y!�DL�/|�El��8���7��t�'?����L X1zb<30�=:\g��:��,���`�i���iq)�`��=�@z�c&�gH�s�ʢ�f�Ԩ^��S��2���/�7�c
O�l1'(!��[��\� @K�����o3��6ꍚ��µ`�0.�1� �p�_4�>M���`��nP��Ju�lWM�l�����cY�(�l��Ak@��Nj7��L;R��	/��#.97}盇��b8"'L��Ȼ��>�id���ɧ\�Vz��_����� ,� ��9zaT�GT���i�/ǰ�+��`!T��4�G��	hƏ1��p!؅���0��lХ|��0��۱�^�w��~���(a�;��$#�����N!β禠��1�����fq��Pο��o.�9���hX7���-�F�6;�L�\z0��%�N]�_� ��f�z���{q*蘆zrv������C�YZ�1a�VRIo]�L�aEU�V�a"�D}��1M*c���<��s�n����-O��'���p\�HP��{�~ ^��^�xCf`�J��LMu�L�>�m��舭��� ��֔���r"�=��g=�n)Rz��l+�3��O/~�u��dl�I�|�h�
o��TI�k�Kq�:F��G��!�}��^{m��AU�O}j�p]]:}��Ma$�%�C�s^/��'�8@��%�N.���oi��#(�93����ц<��?���{�t�ŗ,�?�V�Šk8q"3	���X;����Iq�1�,nM6��mq�G>�ѓΨ&{�zhL�ed�X�|����W����ͦ��}LZ\>�fڳi�t�T%ܝ<�*#\�3��2�*6�g�[�%��1b�A
&2��&d�ɞNT'�zz<������T"����d��O�C ��������@4VG/S G�!�Vw�aql6�}�dqN��kV��5�� vӆ�T�ek��Z���'y��3�`�V��g\�Ĵ�ey}��3�<���#ŧ�����������I}���-0��V�@y���EE2��&�s���֞����#5���������;�#�ӯ~�u�6�p�����Ύ��^&�jeG����z��/|I�ǗIȎc�"��.8DU����ތ���G>RحF#�TY���/:����4YX��D���v�)-�.����%鬳�(�t[���N+˽<A��Օ�0����үQ��l?���80F2��W�i��f-�" �;��/-���)���ۉ�~�w ��5�(��<�����/��,Y/�!kG]vd�����l ��p�
�	�d�l��j<g-r �=�����:hʹR�C����l/��XI{����v��鑏if�r55;Y:Y��n���k��j��ꪸi�o#j�L����!pT��y��5���y�hxv�XHϸ�2.�	}��a�V�Q�~F�ÆŹq��5�Z�C#�X=��L�֘DUU~�3c�gb�`w�ywȆ���*�� �b#���_�bQn�� ���7t3�~���L8���Q�Ϣ6魎E�n-�����ay.e��a��׿����oڃ<1��مt��y@gw�!���n���+nzD�u�U���PoV���{��aA0A�ie�Q|*�������7��9�\�C"�N7�	�>��O;���w��2F���	b/�k�˭���K��3�p`�Jr���Ƴ���1�[/^f��.9�˔�fb��X��E������' X&AA�eʅ�f�`6[���0K����3�%U�#�����|��Ԟٗ��=P�� -�ߝV{˕zb�Ve<��^!46|�� I�6!0�������4�K�����
!Τ�%�i)CCntd\�_^0p���w�l�������k���qI�CU��7*��X����0꾜:��a�kW�zе���"��q����%ȸ���E����X7���a$ ��濺1���Ci~���*��O���Jlj�˱�i��Rߣ�����Eo@Ft=�FٝhηXbD㿑��N]�y"��^Ի�7���=�O�`gp���@���FBc-���%`	%����u��ArU�l�w�u�T��F:�z;�t�x���D��{����Ꙇ�� �p0�ڙ�\���ff| ��MeW� �������6`�N��7���FĜ���&��aM:��T�5�$�[p ��CUi��O��ԙ��E��������9O8d�\�v!>�3���[&��&�| Ev�<t��%�D��u���ۛ�PT�3 �;��z��q��p4�}�����O��9��Q��=�A9��ü�������
�x�\ԑ]2	g���Dܮ��j$���cܙsQ�|:Z]']7ј�z�0�!"V��l��74�&4#�8�u�� ����%��M窚EI����>��-�G�>��^cl:Yg��]ψ��TUmW{���3��Ŵrt��9X���_��-��/s�V�L$'$���� ����-�;�o6s@���(�<1(E�� �IA)Ƅ<��qyŠ��n�Q�9��G'L�j⍳菂�����swpM�nn��6�T����h�h�����u:��	�P��j\D��������i%���l��#�9��V�$q�lU��A�\1�������4`����i1
�D|��jaEN�4�o4���K��<�Ws1_�����orQ}�C�S�+�3ݫT���<��=�C��=!y��6##�p5�O����I&4�yu���J��ʌuZy]f������R�]��vJ�!g����J#��-���'�U��>T�#TI��FP�n�5͋F_�hߊs=[O�m�;���h��n��\��ϢU���-.$���4�n�.78�fLL;�D��5T�pK�/��u��,B��H���^�5O�cu�-�5n���n�R�c)���?=�nէ���P���;�
�űӛ�;�ft���m��H4�,Vw2��vԅ��Z�Z���)��1��(�,��*{N^��#���6d���F��:��sˈ���gh�����k�K�]rNڳ{��Cbڝ=xg�Ӯ�*�{�y�T�k��g.�������ّ��b���t;�y%�?ٱ��J�FqN���ʃ��{�T6���|�M1MuSh��	��`T�6֘Ҵ���\����J,�W�u}�h��u���&������G���E=\��h)=��'��g��r�;��sF��H���?�n�-R@��xs��19�9#d�Nds}hMvb���vYpl^C� ��wJ�q"��!���4ؔ4~q_|f�\��F�ׄ��t�ENc� . -���2Gn[ �ngQ]ǵP��ր	��@aY�(��&6��uy%��e���=���k�s�{u�(ޞٓV��t<3�]{2;���\���SXtņGE_K~�z0�FW�W��r�(J]p���TM���)��,�.�Ӣ�'��t�@����Iw�N�G}��wu�R���Y@]����ˤ�R���kO���0H� &���Iˋ���=,�<)�ͦ��F:|��#��w��f���VTaT��R�A���ޢ+�(7MdU��i��3T4�L;��]���玢*M 0o�^9,t�$��F��u�ܵx'`��ݤ?S�ZA�y��#�ٺ!a��/�fߨ������G�5�]��/�^�)kp�Vj��_����)�0����J:��FqUC3�j�O�+�t������L�=���cX���5�)��Q�ZR�8���������M�c��c%xu�1�6�Y���{-7��MAx��M��z�3�)n_щ^qJ�(]�Q�'{|/��3���Ȥ�P;�	��J�k�K��>��򦏦K/۟���G���۝Ť����®�<��lK������i�I�PWO�uc���i��Ӫ	�Of(�>O�q�~u���z2p|�ȯޅp����`�F��o����� �!�%�3_>l�	U!���u��X�����6"�h��k����:Y*kfiq)}��_I����ӓ���t��Jǎf��ٕ�-��(����-^��Z}�~ҝ/�O�F�C�_�?�Ҳ�$V�u7ʺ5F;�T����n�:����RS��-��Y�hQ�R���5�s�~~~�e�^;2��ǧ���Z�TϏ�i������t���7қ���~�.�g�yR�������Faヰ	�~$���|V7C�� ��d4ҝ����`@k��D���TtC�'{O�5"��m�2��$ǉ���A��n"��`%�B\;4Y6�|��*�~�<�$̣!��;TlH0������'kl2y�`�:��bجW���g��+�7������}��ON睷7u��|;����'�Z�*׮䫞s$�����9�;��ű��N�w���:j�5rwJ�~S���(ߘ\b|�k�_q�h���q�(Fx�'��,������_��1�zu�s)�=�O�<I�����&=�W��>��%���2�Gg|���Q��x4���N8Z��i��t�<W��  f���������<��w���Qw͹�zy-�g�C��Z�ܒD���Moð���)F� �sN��P�{�X�ي��:eذ�]"Q����Xj�Y9���Ψ$jG�<r�h���8�Z��v/��V�3ж��LN�G��z)j'��>C�=U<��umu�`���D����'8�q<tџ4�Tf|0;!VM��1�Zd�3{��^p��:u��|b�M�RUy��,�u[閿�3-/Qv&�R�S�=Wr#�$��I��Q��Pn����H����.q'T�m;�[�,شE��N�s�r�df7u��j9ݩ`�օ�� f���� ��c����9A��djzr�⼀7��]Y-/Z]=8MT��o�RN=zdt2;˼��b��Iw�u_&7�t�E�|+�ػoWQS�
��-k��N�7Zw�mbE�k�q�k�uf<V7��)��MA��sv�dQ�ڼM��`"�	±	�u����ؚ�q�E����w�-�r����R��f暙)�"��ԙ���"���3,Lx<l�ᜰ��u?tq4�E��rӌ��p;-2���9��4�Lk�C-�պ�wBg��׼�ll]r�����a���	C����bXSg�a�k�� �a�a�oX��Du��wDɡ�`�@%�kZ�����Un�Ʒ�$ٮ�g��m G@���5O��y-�:?(�H�Cz�fk��+�̠1>�f4u��ApZ��>#�����ql$�Q]�mLQ��e4K���l�gQ��-�.*�xg����c���n}���3�����T�k��,#���3��52��}/�ڛ!x���K�����t���ґ��y�P�1�q�[o���w{�b��v� W�nd�Vգ�h\U]��X�!l�EU�j2ϭ�D\n(�\#�ȑ`a[+`����9 W�lh.�h����P{L�8+��p�>�&��I�F?�Ra�|+��g�s�>�wϥ�_��t�p73�R�����JZ��`<[�ёw�0��cp��r3 ���g7��X#1���љQ��wx*lxsn������	�t�2Y�����|ŉT_Q\����Z�U�#G����]�RG��ܮaz�k_�.�p&]��+������r�s#ZM�/�r�4O�S,)��������� �e�i5Ĵ{��	6�	ڨqO���QԮ���4���zO�> K�Q}Q�����OY����wo�(Po�$K�?�b �k�G���f���Ͽ�{_I�����������lvP���ٚ�l�\��4���>����>'}�w����URY���-��J.��z����]�˳ҷ�	�9��a�
�p=.^�q���MAx8h�0��0�:�x1)�Ư��x���6M�+�C�k���D.ӌtu ���E�;�^��̦��ܚ�7�^8�Ծ�$*q2ڗ�7TK�>��|�l������C��h]7L�	]d�&Y����4釶���ʄy�f���}�<��l�uт.�#ޏs��PQIX)C�<���Vu�=�#�9�I/%}���h�,}1�2&6[5���n����O��s��tB>_|zgJƲ�\�����ݕ����Һ���:�J��]y�<��oN���E���$��.}�O2��\�`x�x��޴K�an&�(�`7�N��5"EG��O���/�[��t�f�0���AT"��٠l����h^O|��5�\S�g�'�(͝�&��*<͐T����~�+_O���L�+���);�K�~����6*�\)�R�yTÛ�M&,�g��o������IFK���͌s�xND�y"M/1�Ĭ��ɫb"��PĔ�Y������`�(���d7&׻�K�{%F��K�ϴ�i3���6�^&+�O��̂WZyø'}�K�ʠ|����p.�ʹ�{��t��invO��-���8^��h;����������I�Y���s2���<�a�)�S��-t�Pr�.+!���j�<��^z��W��{Τ�9�2LE+�3������:M7�tS9>:��>c�����/y�����t�UW����-��9d����o/;M�B��}|�����A���[I����Z��Z,9���y"��Nǎ؄��@�DZ�Vs.�0e��P���x�p�er4� A��^�<�����9����Lr��i3�>��O;6��Ģ�3�+ L_@4��i�\� g�,��E�K��G03�}��v��Jȵ�t����B��R�'
Õ��c�(j�Z	�ڿ!`��"ޗ�8�_��{���tÇ>��A��I�wq��OJ��|)������)��:I�d���70���^���� %%�ԛ;M�M	��4�~��+��#8w�7g k0��G�Z�CI$��<-�Q{�h5[�����)�1��,�'�ܓӳ�y]ڳg_��ٱa�N&��x �EN:�T��V�K��V]�j��ԔBd�?���.ߛX<V��X�1od���|�]��d�{h�Ҿ����f�f`����nx46$4�9XmuD�iup3�D�&��n'\��O�\UCXN����t�M�T�V@��  ,N6ve��*ki{uۀ  ���+nz�����Zt�����PE=�6K�����Ozz0��O�ռn��u�Z�MGC��s��u[fó��S�Y�UW�K�Kl-�{�/fD�oc�SQ9V��&�8S\�����7JV�x�3������k�9&����=8l�l����+�O5 ƚ��5��d�A�6>���yIf�ץ����j�h;1L@����`�щTL%3�ᛑ-��#�9���`>N\��h� �3�peۃt�H��bR^L��2��8��9�x$�#L�1�-7�J�<`�n����n�r�	
�7bB%��E)�%�j�ZQL��+{�0����^��Έ�6a���(�\�����8ǔ���0������?��-",�Ρ8m��lR�W=��'���[�HEs��H�����3N��B'��%��WRZ.��о�v�=#8X�a/-����[�y���+éj'��-�K���������x�;J?�[���CC�M�o�q�4jL@L"�9�U�P�tp~3F`�VQ8�͕�v��d���i �����~#?��t�W���~=���3�;Zyo��I�P��s��-�Z!��>�/y�K�w��Ǽ�u�+���b'�X��0�z�	�$�LN�����GfJ�~��-<����S+l���TJ�4LH
>�A8�t���I�	u�y�K�9D{栬PF㦿�0M�\��y^�E����cX��0�EC4��ҏ��wu�y�GI��晽v�H�k�Ɏ$��௚�r_���V�r$]x����F�T����.ܥ��<&u����/�{������ )�fc�!K;}�ӟ.����P3��1�>�&��� 5�;*��1:ڊ"��g�������1c���}n2��N���h0��/�,t�W����)`�t*`�e��{'+��Э��2QM�����:)asF�=�O}�:Jv�v�Xz��H���I���4�����ݝ���/�Gjj�	��!J�V���|����{؉T3>��殺���et��Ǩ�nX�fF���h�Z 0aĬ�]�ۚW���7K�RSVE7W��Ut�C��)1'�a��sG76��Dl��Z	�5�܉��s��RF�f�iv�\z�/�<����N��^1|�;s��qX�\j7����uG+�_���n�ES�B5�A�1}�я~��R� ��RmK�q��� ��
��>�s�^�(fx���3
 �G�h���X%qzK����R��L������!|��a1 vI� 8�BG;���� ��yk��s�k�oD������_ˠ����[�^L�������<@�i+���{�&��K���RvTJ��Gm ����H �0�y� �9����3�h,66]Æc����s�噙��!��t�YG�M��:\�M~���]�Q"�𞱁]z,��F!H�w��r�2��N����]��^<v��/9��~B�������L:v,K2�nI�ngf��R��y��ݔ&�rm��7 Q�#ρ�FX�)��4�0�h3�����
=�/��➼4�2���ê�X��;τ�VAv��^p�y�#��~XtK�nR<�)�5�#D�B=1��,s>����ꜛE�e���zX)_��W���J�]�1@#����X1��=������\zFz�k^�f��<p�8_��I�L�s��@nϰ���EO��&[cc>���U%�x3���0K�u?�m���h�tB�l��>�����@+; s�z��u#d�3���"F®)��ҪM�T��y�7��Bj5��K��0�/9��I��,5馛>�>�gQ��ЏN�3����?���l�uE!b��}G��׿��E%A?��.�U</�y�w��]�>%%<�x�3 �/�P�Mi���Ҷ��8��q�]C(��
Z��q�y�s�����bqgh��}��W�� ��Ibuc��T��xH�-����B���qC{�k_[vA���t��t�;���"��qq���2�.��#�/��>������;����oo-�r���L�1�e���"��DܿO��Qׇ���ԍ�X��X����I�J�,�t=&;�`�Sl�ޢ��{B�C2�'��em1��x����~�1�&M���;�K�X�a��fܞ��z��L��+����=���_~�3����ҡ�{�7��t��{K��fs6���R�3>-����y0ȿ�e/+��.��oxCynt�|nE��!�XHb�b1(��(�sn�EyN�Gm�=�G������ڈ���UG4Z�ҵ�[%x����$���ۀ�$oc-��;��+�1������"�y�~����������芟��g��e�q������¤�sh����ӝ?�7}�O�:��U�K�>��H�b�+j�F����Uʲ�Fy�7i�Ֆ�"��XMs�[��m*)���&���b�N���&�Ci�~ΓY�^G�k�s�qm� '�I£
�{9���K��;2��
�3�%�Xa���`�,q}��XŢ=Eo	����õ$@T�"�a�;��owf�sdm��U�������t�������aw�u�T�f��3c�W�,�	(�̪��G�e��������˛���"��;�,+��������x	YS��O�~�����S��k�2H4�L���8����'=��PG�G�V���ʺ]6]���k�ݍ��S��dwٲ�_d
ՀV:a:#�C��ab���\^ӿ�ɕ돆ie9�C?�/��<IF��[�H�_p^>���� =��\�u�-���+�? � �Rg�?���.̦?�fA�U��L��۽׺��k1_�/�L#�� ���h��4�kØ�7���r�fk~Ƞ�E�,��^�}��Q�,[Vա�� A��D�M�!l��WW��J�b���]E���݇Ұ?���ޔe�|��������\e������7� �w�H�آ�J@����'��5�)nk "�D��^�)�|3zOhP��^��	)1���UQJ�4Wv���R�hT��/4\cavRw�f-��."ѰJv삈I5h�υb�c_�җ�����I7�pC�\X0j
\G���?���"]�y�oa~&���H�>��tɥ���fz��}�J���+m�����yo�F�>�g�����:ӭn� .8�n@�ewd0��E&b��9�ew;´�[��
���Pώ�z�-��c�y�v�q|�<,�A��xǄT�SC��W~�p���O�_r@iD_�6Qݻ�s��\u��<R�k�Է'23l�Rg��.zę閯ݟ�C��WJD*�#7e�Z�̂���~��9�x�$���7��<�9�?���T�A�~���wxWi�:q7>]cـb��8~q����X�X���W̭���l�s;��h��y��r*f�|��z����;o�ܰ��sx�)ylԁY"����������$5y5l�I��|�3�)��23Fm	LS��ưL�QZI������_|Af�g�W�+CIU�QXq����vU�S@$~�ӞA&<���T��fM���YwK�Qb�m̱���T�a���*�#�ى��F�I ]�̀  �� @��)1���[�.�c��!��ڊ��kK�aT�`��QEp?H�lJ��j����!�W���if���ϥW����;ߺ?9�/u纽ci�ފU.-/�
+V9\��+V;���'�X՗����o�v�P�oHƀ��싸�}x=n4���x*�4�����}�mu�E�b�*�&/v��@͙�+
Ɇe���Z����g1�E�gXA�F��D�<�'�����u�G}w���)�Y<������t�#���_qQ&�t�b�U���**��J/�~�f��6��D�u�0�L�M�)����n\��N�im��4����U�O��{���(��J��!q|��z�H}.�D�DI�s�o�g���Q��X-id��2�<n�[��/�a�f�XmF�6F���C� ) 0��	k*��}�������e�|.�������͡�OOzʣҿ������Ng�ufa�Ԥ�u�a�_ȼ��p�IG�z^?~�����/�R�PF5>plԑ��Dn��TS���Iċ��Qu�����d�����}#3��p0� ��A����shb�b�1�4�ޱS�!�L�Cǘ�'2X�75�:6un����uT�E��;*�|~�0]}���}�.���X��Υ���i��?-�3#u����q���6N�=c��:˵�.�N����f�Fu��'{�h�ޮ:��D�`��+�v����國sW�<@�8�0b�)`k�M��vp���ͺ@#ܭ`aVW�	���_e���fL�!�s��@o[�_T����iFs��������˳s�t�Ż�Y�^�n���L�qSg&ϙ6*�n��y-���R��0�=��O��C�����Pb��sLc���8�Ք�ԙ�;��6��&��W���y�Z��E�q@����m���F�v���0��i/z����+�t���ID7�>Fk����/f�ѱ��7����Y��q7�9\��E� ��� δ���}���T�$:gG�����A������-}�;�����M3s��޻���eί���/����ԊZ��@�iQ���+����K{�n4.x\`������������4p����:�Ό��.m���ν�U_��A2�Q��	��L�f#�dmH� ����Ju����m.c��8,�kFC]TM߀6b���y��3��D��k^߼��t�_|=�gKY�Ngwcj8��Rf/--Ri��:YR����fSM�S�+=����ځ8��~d�yғ�Tp�M�d`�Ȍ���Ȳ������r�ʪR��$��Ҋ�B 	#$�	!�1k;lf�D���3቙��n�{"�1�&�=xŋڣ��2b�X�&�RH�U�de���߹����n��r�L$���Ro��9��?��1�DԲ�1A��zL��Jrw-�asc��T��v4�[et��)1,�D`�+�ޢ�۽`�{��Ŏ�������Wy����L@���F�dI(�tg��}��Q�#����
�ӟ�L{��L��¿�@�8��}���h����/3w�Y;rx�*���E�;��7��Zb�]���s��(5����yc�6!��� ��Vmh���ă�V�B�K o.���}��7v]S�y,iF��3G�$(.��LR��浤DU�`�(E*�6��������w��W���wJ����pkAj\�}���K����LP���-��_ ����	ϡ���ȋI��趕3Yx@pUL�����?�~#��/�R��ؐ��y�5�p#E���g�
0��_G�)���ø"���F�cUdֻ&�u�N��N�2<�Z��؅0������;Pc��i�3qxϮ)[�De�(�D&U��N�k!�q=�0�J��@�
��#��2����[>��:'¦�C�?��V �r��ӧ���O�f�`�Y�\	s\����K��f�5�d�^?�@=HϹ�+��_�^��u�RE��T��4��ȧ�	ӭy�C��km(\
D=��m��@�����,��Ԥ����"� #n?��|�"���"�6�÷��.���3sԢ�N;�jVo��|���frpWm���|�*�}aN�D{K7���+�^��\W�\��j#a�������g��0b66��J��ؾ�D<�P������g��+:��W�͠7���8���ګ#"��$fg���ِ�'�z)B��'í�!�K���L�Ag��@���X�M^I/X��r7RzLO���&� �$@��85�OڲU�jV_���#ǭ:1c�V�z��v��@�2�IA��D��p�C�\�QQ���8J<��_K��:��ꈥ����leD�����d�S��S��B��Q�{��ET/���6�ݻ0-#� ��}bڎ?a����rXS��%o�	��'S(�j��i�c���*:��a�b~��T?ZK��BlvHҤ��qc�C��y\�{�H��s �T���O�6�|<W=��
�ЩY60�sQ��N��k,��(ّ�XE~u�
t�F3�`���X�Y]�^�Ʌ���|gO�-'v"j���:�!��e/pK�u�7K�L��'���UJa'���!ڝ��}�f6��Õ�9;���?��#�:\m>E �6��>J_��+�����J��L�Z3^�/0՟���|//-��x� ��Bja�.�>�l�Y8%��|���eo?�n��%v���5�#z� �Y�I�)
@'P� v#��<Y�|`�����/��{�Tr�
9 U(2�-!0|�Y
���RܗvQU��<P�XC����W֨v�$�^���I{:�r���ZqY1B"Z��>�������_�'q��\�zΐ��@�K���޲\B޻ m��@����]��a�hu欓�;x�����_{o��ɤƦ0�[Mc}�,:h5$jM$����������a����К�R	m ���rΫ�._�����z��h��>�e܉�O[��`�j�6o�loy�+�U��>��k3��T�@��Y��rS~r�z+%�2f��e��sA���u��l��7�
����=@����x�8"��:Nc��2/D�����*�ʟ�&F(��,�m�\o�s�O �Nf��Z�bZN�t�dgR�W����A��%��x�(�׏ϸ��`�Y����Oy�=�'Æ7|��1	b�FY�];��J�c�d�S[�f3�n���[��軒Յ.{#�!Gq1�!|���a!?^�"����(�96h<�~	x�3�j5��rA���m�<k5�X�����42����~K�[l߾zn �t��@_c�&�����20{젚��^T��� �0	���SQ	�U=t�✹&@�Ď�^AJ�i]�������~
�N'�\��70�-��kWzX�ۄd`P#�������yp�� RM����T%x���lI�A��B�n������l�[n�:습���v���WZ��l�&vx5���݇��Q�<?��w��Q4�h��9y��=s�{�]��=AF%��ǺQJ��0�[aݶ�6Q��q�ngE�x����W��]q�Kl�maΕ�L� uv[�Z.j>�G��(�P̛����9W�DEo�(F[ ���q�W�e,S�>����6Y�`/�&]7l���p����jt����A��~/ZD�����-��	<|��>�Ĉa�P�E�����}Z���[��'�x���w�զ'7[�r4�6�<l9��WJE� M4���\�0���?�/��V<�sL�gi�Ӧx*�ޜ�?�Mb9 X��d{3"�z��A��Bs{�d�)��v5��i�����J��r����ޯ��/�gs���_�2H��1�p30s��Mo��n����&)�3!^U�DEb"���H/=��5ߕU���1�:����=��/�^�#!�ƒ�-2�Ҟx���GK��r>�8A�*�����Jr����b`� �{
�}���&s<�[�m[w�S=i��������ο��p�J�̇�N���CE.�G�y#���'�7��P1<�/B����s��h��o�ɴ�EYW�zf�(�X ���"������e2es-�]T��̘� `��>��v`���n='���/b��S]R6�����^۽߭�Z�&5�"D闯�&WL�_ᑷ5q�2���^Hܸ���=�y�s7�k�.U�>މ7��jJ$�7�sG~��8�;�{=�����Hw�c*��E]�o�~ǿ�ı�yX2e�����_&I5`������ӵ~ވ�j��J���@9��I��z�i�������$�C1��O�q��j�<W/	�or�7�&��U��B/���@�Y�7h�o��"�� .h�X�_t_������'҂�����W�)�iX��\fv�ZSv]�*Q�011�3X��^hԛ��Oe* �YX��ʞ�d��_�
@��4wG1"а�?����������=��Q9Y�U1��I~2�z�Bq-���������/��}8퉙8�ʕ�.��۹k{xo��t��V�~}9��"�<�]�[�=��O~qkg����{ ��{Bxg-t/�d��-N�a�i?a�!Ë�:��j)��_ۻ�s�ħ�/�G?���`T�t���W1^��g染�,λ#zfE��v����E���Q7�'a��}�;��Fy��/8���^��:1��j�
�����[�;�EXj�+���Qs�8��ڄ<���or�I����,pdE.�����Z�IEU������{&�ũ=}�i;}�6{�O���\p���(���u%�ig�o���2�[��" V[��P��s�꓀ƃ��"�i<}ٖa��Un�=��Kaq��f��C�ߨ��B��p����"��9�9�^>�gy��1}���W�U{�$��o vo��QHs�?{?��}nkKX�[1,���6��6��j?��[��~hG�խ�:fI�a�f%��$�eU����W��=ޟ7L�YOZ�\�߰�S��r�=jw�R�k��5�c�up�����;��sv�%[�y/8;L��(&MLe��-���p�J��(2���U\�9��yqT���X/���_��׵�3�F3��},r��V5>BI�F��g
�;/m	��o��R'���6z�H/�K��P ��`��I��W�����"�΢$�LR��jiZ�� '� 5�L���y��߿~������y{Ίf�y�! �i� ���)�Zq�x�f�r�.5Ǉm��1�QHcA��rF2��-�P�IQ��5���S�m�z?Q�����v�i��~��sΌ9�X�[���U�����Y;v4tvi,	�X����٢�������@�"Ǩ1й�ĮS�D�g���^>ۛ^���{q3� z^-N�Q.I�|tm���;���{�aݛ�DG������˟�!xc�f��]	g��� u�R�)SB��n\/�2��Пٖ ƍ�V�{ٕvڶ���ө9J�g#�q�,J��d�5���Z\�K6���AK�?�v���%#�hʸc��R��*Z�}���P���z}�?����そ-�,J��a�}�DԋA�*ۉO�7��7�f�UȎ��r|M��e'�fƾ=ŅU����1g4+��8*n
zv��w��O��^* q��+��7ho����?k]S����(��{5Ű>�;Iҵ�;IR#�;^}��QR��&�$!���VQa~�VL_����[�,��=��>�����֌I�[��"�N��ju�QNia!l�]���������_��r�Z���.ُt0��r�=��T<]!��NfolO$~�{����b'�J��|������|��B\U�J$C9f��sv`5��Rn�"�S���}<�P�,+��Pa��E����K_����}���A��V䊼�<g\��.W�T_4��,j�{�N.WV*ZI�>
|�a�f�5���>A")r�(ɍ�L�GD��z8��TT�����&�K��J���I4(�����s?r��ү� Ҫ���)t�k���A��aR]�y?Ӫ�����X���i�gp��⮏؇>�ak��Z�bڦ�7�UW���\p�5[��)�5�>�w�D�a�����U��8�Y1LE��4�+�%G +�b�_2y��{Y��QT}�W/����@�pjo���!����ჶ0Oٓ�0qjv����z��l��C��o^I �e�n��D��$�E}��d���s���< �L��b�J�_��m����< �"� P ��r����W���=�^ �$D� ��|~��⺤?����??r�@�������ƈ���8s�~ ��e�+�\� K}�Ky����RO �ܟc g�!<�M�~��D���򒍣����D���&lQ�09U�Ns��	\/Z̪5IY�mZ����=}��0U*fn<ƭ�s�Ԧ�S3n�8R���o� �MP�N��J(]%j��	N8)����pd]O��"�V%d/�	KnT��0�8e���l� Z�<���x�x p#*�B�#�|)}�>H�H�I�3�Q(Iw�1 �<����v�B�bY� �!���$} �'�61�C�u�^K� �~��u���.5цqEu�(Ւ6C�K^���o�̓��92'8_9 ������w�7%�`���"�2/�@"���k"��]f��}+�������L0�h#��h#���+���6����?ǒ��{r,� �	k�{2wi3k��Tƞ́$2 k�q�����_�r{
������w|j4~����uJ��a�F7ϰ�5լ�ZxtSd��j��kA
	��MQ�#KE���'�c"��j�y5�E����E~���}}���>� �+U$�}�+l���)V��><#ի��t��X�u;��p,;==K�3Q�<I�(&��_n�^zi��|k��`�3AI/�����n׿�;"xS��s�+��"r=>�`�Dz@��E/z�IA�J�mǎ�0��m��CN�(�M�O����7��3�ѵ~*˥��W��O�FLyOx=����|_�qC�TE@/�CWCE���g
�3��c����U�u�ߜ�Q�X�w1��1?�r`�q?�x����[����7P����CF=y+(_,m%/�R�z��P�[ 5�q]@S��5�Us���b� �!�2����e�P��,�	��)R�E����l�36���X�h"�&lێ-��+/����\km�=�0��Jo̕��3	��gI��T�����͑�����G�#�LT���K6=*� }�I{���:TL��Vj3~�G��E��讽N�RIڝ�M���'����n��^xQ �kbZ80�k�d�<&���&zB�DDB&c��B�g�g#�������}Q�p�7F �a ��\�EḰ�� <Q��^����D%�Ī��Q%��������3����
���Im��~�?���N�YXԅ�[�i�86J�Q<�$=x��]!�S�aj&�=�L���	�c�Ј�,0/��V��H t�|f����8�9(�8�y�F�25�#��1��X��E*#�a��\-t����VF/Iq�Q���y�C<�r�;�t��}���Q��aé�r���2��܉#�%aOڵ];�����F��/��Z���0��Mx�V�Z�6=#�2�[����I��V�4&��+^�
���ۣ�8�ӗ���1/0e��z��C������|��:,���4���x���Y�<�����v��),a��M�,�Ns�n>�l^t��t��ag:�W�
΀�!�p`�Ʌ�]���j�}�����ʎ��"c����Q��w�i?��?o�''+��u��H�-��h�����ݴ�w�<,���/>m�f��E�jŹ�>�F=p�)���֫5�u�^U�d4!5h����NznΨ�5�����,nE���s�3��� ̢�w�ׇ"�|q&޸��<wDI�f��X�,�é>`�����.d^�^|Fg�x����u��F_�I��SqJ�bh �J��A�h?��E����0�6m� �\�)��?sԵٙ �NV���F�c�[&�3�Zu"H*iۦj����M+U��Z��e`�ݾ;$�P�UkC���������+_���9�o|�#C���I�>��&ȳG�T��넥�{�,��!�0�G ��Z)�px�k�	��(6��M�͛���l�� ؝��yf���	�>ɧ�I�?X{:���.�"���R u�kq>0"����ܱv1_tO�$��7t9G�Өpן��sׄ���l��M��Hy�p�q�y�r"�[=��N��0#����H-�QRzMMl�V�<�Oj�0���a@�O�(�PŰk��7@���b��es�).�k�P9��ec���9ǵ8���5�
��\����yϢ��zp���,\��p�p�������%��}�o='����0�5N~��S�	j4�1Z7m���
���4�ԷT����߶˞s��>繡�%�Q�+�$�����_�U�!�C����s�p�s��%%�o��Jq<c+@FR�馛�3a��5�^�%FI�<�c޾�/������/�g(}�����%��������&���9�X�ͯ?d���ý^�`Lnu��G�k��6.�,nC��{<�������|�#��?��?�7����Ap�StA�`�]����:e��_~�����oٿ��_�߷r���|4ט(���4L� @�B,�|�m�5�G��a<�4P7�:r	[�3�rh�J��\@J�x� ��yϕ�����g�J���E`�$��F��@��a� �Ap�0��o�}��ĸs���}U�$�F	�̱0J 8�7��b��pq\��dh�I�+ΐ�2��8�L*>֟�����$L"�N�n�#�Gn�F����������{���j�˿��&'�m���"��������$�Vyn��u��W��mx����'���}�8Tm�b�Ĥ��c�d^������u��'H�K�bs��{����VXop�k�����Q��������"b�1�i�2�h��XJ�"]��3vFO��f��Q���ɋ�C�̄G��7��w<����"��t�ϖ��M�y�t���#v�'ﵟ|�+���P9n*����fä�M�Vޏ뽎S�n-4�>7,���=�z�azY��E ^Kf8ԟ$�le�l�SD<t��@%zz�"�1�Ƙ,��A�����\��z衞�!b��ay!��l	�7��g�T 9��& * G���Gnm*���K��fA������c��J�����s���稛�Ƶ��n+z�;ٸ;ڱO}�s�������4+'�Y���l�1�5b����?��`l��/��^��WG	��t�a�P�s�=��s57 l �b~@|���֐rxh��yހ�7�7U��P����a�	H�ؑy2LT'�.�{�!��3���#��YF&;��/t�I̎�N�D�a` �{����4zd:����_��x.��E��̊�;>�x�ĂQ(v�DÞzr�]tɥF��VNx2���Rf�[f�r��񐨥�#ø�a���)�P�/��$2�3�@~���R�9 ��� Wɜ�h"j	���3��׼xj�h5�2h�!	�4�>_5s�{���7�q�=��I�r���K�"-|��w|���*�#��!{�|���q��~��:>P�$�>E2�J�)1?6����$fJK����
���u�)�I�կ��??/�O�������8Ό��-�_lzR�ȷXz[ ��Fg�f���o0~y5�X�3|V�E�2w��
a�k�	'�r�M��	�X�t+t�"�GG�k�B)�(�Cް^'H(����u������-�qD8�l�z
0���s�uH���=�)����6�NY)�����n{.:7�T��V�\�ʢ��tn.�D=��* ����`H��wYS;�G��-F���������~�^�Q�;�"�2X�T= �`?�R%� MZ�s�������@T�u����	�5�l�"����B  u��@�W��j-x ѫ���ŤDޯU�О��5�s뙣0��N��ȅ0|[� �i&�����OX'��|c. ��L[XC�6y��ܐ��m���*�:yI<I�P�T$�1��JqTr��v#y��j����ل����J���	C�i���k��хl��YR��N�T4��Kc�2h�J8!������G���:�� j�c��B k�ypF�R+�F��sv؏���p�r����=�U�������D7j{1�b�������yė@g�ܚ���3+�L�mY)yN��?f��kMî9N
�������N�F�v�bëE`�����^y�=���F�4;|�`�/��.���S���0��,��#�/���XI8Tc�(�$oFa��d�+[æ�C}�6�  ��IDAT�{�jS�����ݼ_N8 �8t9���[e�G2����h�XVj-h݂�ᢆn��[o��	_��1�NZ�F,�.�M�Atmj�do����=n�+_p�M̴�Qϸ�Nhnti�p�#R��'��9*m�E�ٝ%���!�sJ�@U . �$V���=j\�3��Î�z����\�z�0�|Q
7�0����n�C"��+i�!\J�����_�cs�;v��^h_r�=��&gg�n"��U��\�U?��i���} �ԋ0(��N~�#�$8�G��! �^]���$n��:FҔ�^��Ͷ·N��ˣ%�m�5�Һ��G�����@ ��7s����� P@����G��N�k�1�<<)=4�HK��\���E�{l.j��]��l�.6�#v����n��a�L����yu��&�KDU�5�"?Y�ּ�B",˫d��s5 ���Z�"�֥���~����b؞
��u�Q��b��:ܵ%|�����a=LN����a������mێ�;�[ϳ�~�` ް��Sf�w�.y��֩�\�ۆХÄ��o��0���>�v�0e��B>�M82�z�(5�����z�a����n�[.-.�xB��&β�A]�:#�_�ThpQ����������K��p��{�[�b����i��{���g��6�t;�|?���|�R;�[��������a��)|��N�D��FgI#l�$@+���Pz?/�+��(�k\��B���*ǩ��Ѩ�4��1~W���{H��c~��+w��p���@�dڴ90@Uk.�b����}���Y����?�J�6���ێ�B��wZRg���|��	k��s< X��{���{��8E4�ە@@�A.i�� o�	�e��Ƒ��K�Nw��5J�v*=G\i���v��¾3ޥH@Z�pQ��nG�uL�k����aN�~Ǻ�կ~5�������Q�|�3���ǃpֿn����_�;v䐕*d|j9|�m9�:s����Ls�\��H(��,�Ч��n\㢉(5�al���Y>�D���E��ն� <
�W�E�jQ�����b.~�/�� U��%e[�_�|�c������8d��MdJ�b7��j��Tmr*��0g۪��/V�2^r3U�� F\$����ߏyq��-�H�X�!�&x�Q_�ˋiz�K�R22ڥ,o���I��n�V��XQy#�h"��:�E����x7o$�3.':ݢ1�Dˑ�G�O�/L�b���3(ɱ�J}PKc�σ�f�-V�$a"a<(��<��Ӯ�a���9g\BU����ë �,�q��ǥ/�q� %#�Oj����J��aTԉS?�>+1>���j�.v9���j��6�g'�B� NNLe��e�I\A��R5��n�gm����|�N�~��̐U�eR^bY�BI�a���d��F+\�X����C���M .�_p��3C�Ǎ���KF���q������{��R��5�Nڕ�#�����p�sϏb�	�%=O��_��1*@C9\��A�NGu�)K��irD̡�G�Agg$���g�:I���V^?]�K�-P�_��j�H�X��Z����J �ސF���ؤ�ܘ�Ae�řӉj�h��o~�+��-�������)�J�s�Ji�Jf�x����(z���&�Fcr`���F e�%Ҙ����T��~������%i7�7�W��>�ASSS�Q#X�w±pɄ����������~�5a�̎���XT��{W@��9C� �|0Hђ��y��-�(�BZ�M<n<55w"�.����H�� ��=ј�n��%�����̎�O1���:��D�d�#a@��1�	���5n+<��ﾻ��ɷ�{pm�����p�u�f�b��J9��ɔ�����M��C�	�K��W�f%��C"���;��+TG��{*r�Ec�8�wW�T[ƵkԹ�8�����h�x=A�_"�&��e��d�sRH�KO�6��8�G�ݳ1�?W+p��#>}�v�/��?�Z�;�
��l�MK���=�	n��{���Ђ?��?s�p�hH�G�-; �8��+�/8�ڒ�?
��:St�sA"������6���^�F�N��ֆ�$�s��2cO�����^���Fu�SO����>���a���� H �`��JN�Ί~"<��?��?�����ꝏ[�|#dD<�8!];&�ڊUx5�r+�؇��]ĕ� �͘O�r-���������~4�C1N~`t���a���n�=[���V �e�6{�Ͻ�~��o��Z �:�Y�&�a}&��%������E����N�5��;�w3�E-b XA�ɢF�@����%&��j'�va��سgO�d�/� |P�����R���3DFGp��Db�i��^-�	�I�XF��$��:���c�Չ^M7���h,�T�'�T�$r�:y�]��^٬C���[b;%NhW�@��A�c٦&7��][�J;2�ɠ�8�<� .��Vb��aI)��6h�����T�42@m۾c��s޶�VH_9���w����o�s�6Mo�)/QS�N�*62N˾��pq� . ���uWK�T�J�$��WG��^�
��ʵ�����w��3�( ��b�b�Pn�bދ��r"�25��dL�sքƱ���_���z��#Gˀ�FB����B
��X�6�T.��蠀����t�ܓ�Jގ�T��+]��q醉�==k؁��ؾ�����fw���љЯ���m�����a�V�Ֆ���O��A�σ��4�ymCkY�q�&����ڷ��d`��
�q]S�sj����/ ��>S� ��T�p�bʊ�%U�����6@ޣ�p/WO��&Q ��6�?���PR�3,�'V	K����Vo.D�����"G���N�)3(
�``v+v!�F�w�*�Ă��ك���׼�78��2@�Oj�z>�ם��Ժ�m�|�}꣟��O�#?x�����ض�;�`i���M�;��,����l���$��X�� �Z���\îҲ�����7��v�������v���ע��4�b�����Ի�*��u�]9R���J��J����� ļ�������B�;`^!��Yد����Ғ �@�)2��-���H�tsp��P\�"�a��v���9%�� H^9�F��
�O�B ���Q^ �{����6��'�x��򃟴׽�v��=-�GIE8�wx���E� ޠ���D�i*�&ʹ���0>��O��s69qF��b�2x��,�� �:�0惫�//@���4�0�!�D;>�I*	�����&�
?1�ΐ�׆��5�R).��h<�Ԋ�^�8.��U;�>3�Ocu �Vɪ���3�C���2(��b�xQl+����������@. UjA�, JVI��g�*z@���R���V���{roVl�����ٌ	���;Q��A���r���ј��Z��o��������c�nٹ�LS�=�q��R|��ԕ+�{H�VjD�2�B��T`�7��W^	~$|.j>s=��Sp�H��ʹ�
�����.��}n�4��>.u@�\NN,�̦�x��b'f���є�V:9�= [t�@� aY�"qB�t\�xK�C�1��AɿP)� �W�|�'�*�z���|Ĭ6�Yi؅�m;N�l�S��ޯ���)��ōN;����ڠ]DE\cYǋM@2 �T%��-v����_�o�*�^�lW��B��^�1[=&/̏-���*F�J���>�X�J �+^�n�a�|ДWcB*X!X�}r��֞NZ�4�#r�t�U�([ϐ7�@�H�G�x7�������XY6�ex|>
��j������O4��w��t������ُ��z��2ʦ���9�T�F�{��h�c��Sk�:t�<�6��r�>����҉k��X*}^4Lx������#�8����+�Sc���}���?�$-?��w\π?6sIMJE꟭o��->E���[|��L_�NJsHY�._��V{�<�k�0��}r%1!�̫V����*�ʡ 	Q^GR���)l]��x`Z��گs��y�c��� ���o���ਕ���ݑ��LD״ޜL��R�+��杘6�&�<��Q�����1�L ��>�s��Џ�;>Y�`�Rߓ���G9����,��8�-�[@��V� ��xw�!4�p�/;a�N���[�KΰK/=�&�Kv���3S5�cXr߻�%����DrX��F�o-7I��W@L�ߚl���&���姩��r��Z#_j��=�H|���r q���ʷ[�ڐ6I?*䟵 �K>Z��_R�(O�����;��RV�%SH�.}cqS���}qU��6IH̊6X�]I�z>>$]�D�/%5��R����7�{����͛lbj2���\w����
{������3b�#\:kթ�����w�����*Z�&T����
q?��m_iE�C�'�(MWǍ�>�����/山��a	b��<�����	9�m��l��Y|�v��������9�7��2CC�'�.�W[.YV[��J��>���X���.U����xx�b��B�X!��6Gq�R'	�]+$T\�mD ��8�︎rp=y���(N�K;j���|�ө��F_�Sz?-lq��bf.�y�bD�U�C��,����$�{��Ӹ*����K�.���a��E��j�/4cy���b��n�풋ϳ�]fss-k�� Y�H���kw���h�h�9��43��+!yRx�P��J��an�9�F��	�;&{�Cn�}����K����&�v2-�QC�������M��i�Z���>:g[gϲ��<1��sP�#N�W� �}�-V��L�,�Sq�J$.S��D@ ��X�ճD��-p����%���(#վw�����H�Tj3��i��y�R�S-7�kN���j���ࢴ8���(Jn}�(4����^��D�}���o�z�r���m0^#�Z�**È��#���FO�jeҞ�7g_{��<�0�l��B7[703��1��Z����3�Tb<����o��Wh� �dFp�˹�l[?�[A��Q;��Z���RWxqP �wT$5�|�.ngs'�W��v�:h� Tu���g�D�F�'7e�"ba�NLa�Df8/���*	)����������1Y<�Q
Pe'�q��	I|g!(���ŕK� (��W�G "}1�䪦"qO�*ݭ6��A{U ק����p=�)�c�VMqഏkpm~�]��~�-\[ܳ'�M`��Xc+���zR�����1��6L���b(�����p�R6�N��@Kܼ�U̢�^�g�ev�;z���߹�����4�Sj�I;|���}���u7��]gY�4��b<Ƣ�/�8�� ��y߼$뙸�H:����\n�9�xUߊ��'��������M���vs�Њ"?f����>wb��'�:Ĩ01�h���	 ^�n���s������	[?��~� 	���cq�X &�^��^�X�8� *�-w 
�)~�J~����$�^zit�Q�@��K!^/������x~���8�w��{"�����M���{|�rJ۩���'ek�$��]ʅ�爣�t�RPEW�� �#��O��v��2(������n�#��$ƕ��MQ�p1�2���H��u�;!���>JGK�i�*�r�+��N�6	t"��"�h3�*T�gGpנ���2^�햔óճ���I�6�FN��X��^I�U��'m ���{yھ��w�G�.xS�Y�ͨ#�:�#q�^�(R�.?�8�w�%^�9�	\�{�����5��sZn��%�T������u\6�S�5�-kwI��-��0��NసVu*��rFT�]�I�"���ʑJ%j���ű�	�Q��N
P�  ����>�� G\v�����ߜOi�����+��"�/`��v���  ~�>�`�� m!3ɺ �.� Ĺ��`M`��T��K{9�� � �r_Tuc�����f��崝1�ܛό# ��*}.?S� ���r-��f��f$� �6����@9�񑏻���w υsy�<��&b�1�;�:���z�$��� @�b�3�����G����9�TX.%�N��2F-�AR�&Y��tлD�J�3ʯz��焇q�ˡnw��	Ot:�ҞRO��*�x�b����E�U{u�#Y�ДA�u�]�n#N���;t`�@����dح��a�΍p�ˢ�?�<�_�D���Ćdܒ�	�L�Z�3�� �D�X�$,\@���x�c��NΉ�R% . ��� h�� `D;��-�K,.�������m��s.`�m�x��q-H�5zv�E�JWʸ�+���u�I;��6p]ڦ�d�4 j���6 `l!�9%cýd�U\3@�̹\������fD{�� ��OWc���<S�XQ(�TO�������`֓�;b�S5k�p�u�<S��;�0*ktӆ�_��g�c�\}����9���uV�R��D_;�	R�TORE%�Ai��ԁ^R�h�@��ƌ�n�B�wB�b*���muc"5���kAIg'qKzE�(�1�<�(~ �u�� H`��`��y\������9'��J%�햛�cS��z��&j%k5J��ɖ���;��G�Y+��="�Mn���W@�� ��{,�0u�҆�Dn?�;:�K�'�����쾺3�	��BC!�ø3�(s@���9�c/�<+�hh�D%��$��Y�� ����/s�Ϝ�=�N� J��xp> H[�tʊ����q�@��sƐ�܇y�J�|T2���U���O�c�#��VF;qb|��*1���޵�����C� 6>�'����G�.���).	s�����ǣv���so�I{�-W��dhC�n��R�[lrb�-,�y&���	c���G%F�A�#	W�S����|�Oگ�. �������9j�C",��]�*�{ch�9�n))U˕�g9 �lpR,�t���*E�%݊&��E���a�8Y����t�,UP�N��]�;`{�O�=I���~�v۱}6֜�v�V�۬�[���1��s�>aϏ&�����A��Ȋ�o�	q�qg�XIO�o�	 �ɨx{�ѽ!D28�y ��3D)U�P2����K[�r�&��ui��^����W�'O�B�űÙ�8SUX��T9^_�O�6-T&������㽌\���r	 �pќ#��r�p>=���4��kr,��o~����I{�'����b#�06����H9O�gq�P!�v]�)��UJ�5�l��	��bpu�[8f�v��O�N�ԯ�����a���\���V�6D��v�|e���@ء�^̋���xx?t�����P�Yv	��}�Oi�������N�'��.��J��KY�Z�U�?��N��w�]�	�B�=��.���jb�kP09`Y�e ����鑊�vSQ����!;��vÍ�И�a�[�Ul~�p���p�eu�'�·*�_�\�
�3�f�͸*��W�B� ~��+_g<�^g��H���4�p,|~c�s�V��3���(��Z�<x�'�����N\���k�����f�zCB\�<+Tq�X��Q &�����9G�>��NT0R�p�Bh[��8��~P�	`�g�ϱ�j,�K����5.�˜��8*�>�y�kȅϯ�����c��-�a�զ�9n�G�m��?f���vɥׄ��u��Zb�z7��"�$ϙ��|7�օ�Ah���}��T\�gc��O�m�k2y6��4/�!K��p%�N�ֺ�r�SI��ݥ��%I2	M��o?=r  �V�5$�*�c�9�ゃ�k����K,�$�L��0&?�0]��2�(Z�����q-���B���"7�o�-a��ڑ�lfS)<�N�QˀXE=#wrP^? �����&���r�J�˱��G8+���� ��=L*��x&;�	�p<�l���\ �de|y��$�ȆH)��\�x�<s 
�gŽ8O�)8y%a�E{T6_ �v�0����617��ע��ƫjJ���C�i�Wp���h<���W�1��1�<��8T�)�8c+uc�x�,�+m�m|��d�L��T%��gB��ӆ!O�u���~��b�l�X�1�O��b�>����w���֨W�~����v��o����R�<���`�~�T@�� ~�y�KV�"���j<4��K��ld|׫M��y��F��#�e�+r��Zµn'�R�s	�!p����v�,����.�k����)�� ��o�ǔ�c�P���cLbb2�$���K�����U��7p����8pЧ?��\^"�(gu�	�,%��v+�;����vϧ?o�yͭ1�O�Ӵ�MC���:�����[��0F,x9������?�X�Ð�X��])�����(%�:��s#LD&(�v ,�ǳи�:
�г���t˼�N�$��㸮T
����C�^q����7��g@�k�l ���o��y1�|/� s��.��`^z��IZ�pO�Oq��2�%�}%Y�_��I��gmb���U�z�}qf��/~�0s�fd/(��u��U�am���S�Q��ԩ/�����=�������T�t+'ӱ��f�oe%�� K�qw�qG�����!)in���{�9I�+{�|đ� o0HA/�S� �1e�W�B���=7I�2@��T�+�%]�*�0���Xc.�i�p�<Q�s��+k\p�E�E���!
�O�!:&�@
7C� 
�]D�4�p��	1F�ǽH�|�7Dq�kHL�V̆��g��'�\�&O- FXDO<f\tVh5�8eN[_�����~�H��s&()��p�^���s�3�OARoh2KO�݅(p�2�
|� 4һ�;���>�d\��(	��) 7��k'5��?�%N^��?�M�`�'����"����K���2
�~�W�\����MB���`L7qc
~Иs��q�0���$$�D!��j=�:O�M�x"�#+��j�yZ�	�0s;AWO4�-# �Fla�y�k_�����7���_��h$��<|$����{���o����iH0���#�y��`n�����ճ�z�W����{G��J���R�8���-���XE�`�����tǄ��Q���&5�V�X<tL�*E�l &�o��oG���^�:���?��k���o�Piw*& )�L��τ�|�.��t�𢳣:��l���"��,�{&9ur��J?��:�/����o4Y']�<Ε�����k  �X%��\�+xC�S�%�{�I4=�-�M%��.�N�~s����w��T	>���@��~kj��W�s}��tw��i�)��kjQ���8E ���&�!�u-�Qu�I94��q�&�st��W�K�K�ubn>����NEIy��;m��h[1x�"�����Q6�'�O�^ �+�XA�"� E��Cf|��К�3���*<�Z�瞽!�k=��Q�^������C�k���@���ђ�p���X�ʅL�ո��K���1=��
~�|�m��tϋ_��o��A;:�����>f��[��.��!#�w+iaxn��p��mb*v����{���Mw�y�i�a�3�r�R��rN*���YC���3����E��G��G�����=�h�c�}"�aM�H=����x�s�
�+�&?�ݑ��Z�i��%�(oȟ�=n�ʵ����@)/���,JUޖ��R�/N,��J�����a�z���^���I�T>�k=�����,X��h�R5��nD�6���U��;��}v�ȂMLZ��C{�S�c�Uצ^���h�;��^��F�����_��CG�J��ɥ�'�B� ���1>��&�ׄ{����o�b����jkN0!�ݩ5vQ�&jUk/�^�'C7s�aW`p����bO��B�iBH��$B�HG�%�R�����ϸ�� ;��� � 2���}�}�*��g`b&kv�ۛ��v�%����1`��Y��8���'^p��][���o�I�*���Ӱ�x�����N�c��ŰW��W��ڤW�J�H,�P`Qz�ܠw��QM��}_�F�߆����v�����1)��u=��k��|��~�-������^m�c��J�i+��9��*���I���DVmrz��Aj��*�5/��~��������q��m�\���P����f>c�Fs`^+i�ThzN��jozӛ"|��}��2.�%T��n$)�5��M	]�ʪ�,TZ��X��<`�6g�Q�̑)�I�_�.jI���S��4b�2A�β#��t
�I<7��g+w��,ƀ1��Yq�pw�}w�0����-G��܀��D�����Rb[wL�� }��۱#�6�y{x0-�7�<��-�Z醋f}*�AkA���5^I�R
LWg��������T'��vع{���?�Ή��'�mj:K�Z)�֤��b�@�D
�6*OT� ����ƜB�yEj�0:+镘6y�h��+�א���_hp�{t|&��C�F6�iH��j/� ��l�F�L�ð�J=Ile�؉����DW��Y�pź�@��)b���$���x8Oj����%DN;6ޡ��쑇�N��Ѱv�Px�m����ID]���Jv��nu܆���~��l�=[��z	�p���ѣ���=�����*�n��F:�险 IS����K���"y�H�º7b=���+jL_�G��C�k�pˀ/x!5��aĠ'�D��M�eWP�*�,��̛&�%�n
Lv�P���N��ɸ��������4K3X�(S��qH�|Fe��d�fgH�++�z�w��Q1���g�$B`��J���Ur<�B����lM�7�}��k�a�MTÎ����I3�N���eJ�c��X�z�σlэN�A�l�L�6�@{z��������]�G�o��]`�]���%_>���zLeI>a��T#RN�fP
(Y|/?ie��3�AZ��Y��>��0�'=��G��s��K������S�k��hRD�7���+� ��EQ;R_x_\����^~� ��IB�) �?��?���>�яFu�9�3p�8��.���Mo��`f�q��ܿhS;-��lf�|�zb�3a� �M��i+(m4H=\<�67h����nVA���ٰ~�n��Ԍu��ӭL�x��>N��f��J����XC�h���Ry����3:]�{Yìk�<X>��OE��t�rS�a�����e8�1+H���}B~�5ہq��ڃp��q��[7�F1B�R|\6����Y\ ���y�\A��c{�SH�p+y����z�1�@[ ��N+� {p�|��d �f �2b�Bh�p�.�ռ�\��a�;bm�����\?���ؠg7��\�
k(H�ݬ���d��S���歜�����vn�f�o�7��pl�q��rC������;�c��^��UKF}T������䋷A�;�D�3�	�꣇-�R)|^���J�Y���_�L��Q;Yp��w'����+������z�������=��w�;�K_�R{���B�ey�h��So�;�D���$:jIe��{�b,@��'73��#ùS6�诺�q��қ�Rܰo����mг��:���4�`Ǐ��v�F-s��t�T �ik^�%7<�v��8�i���j�u�}�=k��W��r;`��B
�Cc>^Q>�V���E�D�*I[�
k�y���}��T�]-W�n�j����	�y]�#��V;A�6�w��."���h�"����9�o�v-�E���+�J~����?��N��R�U��ꂼ�dR
��> ��ІFhx��l�&'6�wz����-;xpq]�����'��z�S�ݍz� ���Ӧ�mo{���c���I���Z,��l�lz�Lkf�Ըa%�'��T�eyT�
C�o�u"����3�>�$jSHҲ�	�A���w�ԧ�QT:S��@���D�:I��D�Aة#�IT��J�ȳ�y6�GwIE�� �+6���?�{|������y���}�I��
����$����f�mE�h�j2�w6�9۶���0/)����I�C��½&��J2��RF9=<��
1��J�$�J��g�����S�7�'6h�i��N�Bnz�@$��V'���k���g��/<C�1ĵZU{|�U&f������z�b�F�T�6vDӱ���Cs ����f����������/^c�S�#q��-˭<#8߫E�6�^ .�֟v�̱.qW��y���'�H�Ġ��^�je��8"Kv�
�KΉ:٣O�%��Q����X}�+���s W>+K�t5R���!:#`�w��X��F/��"��8�Z�G�_.��L��#����]x��v�M/�͛C��cG�
�KF�0q�R�3�� ��<n��9o��mp�]��'.bra&�c�R�@6 x��i*��;�T�3�1�J˶l��c'��?�����+��Ѷ���`��-�N[y*����n�lO;mG\D�¬��y���ڽ���ɵM���`��d�)Xs>�]�
��L*<���'�e��e0�Y�$O�ߍZ�Ռ�xN�UNcxa�"�~��N�Z�}AVS��а'�Tt�D����1��j�XDՀ:]��#�b�0a������薆h0)q����.�Ї>sI�d<\��[����8�سx\7|�e�t��G?�����7����s�ґX#�رV>Lr�
��˃����76�c�q`d�/�`�qL �q$��mг�2Õſjd��������~�ؓ���W�������R
@�Uo��a�#7�l��������7�9d�(�>p_#�Ǒ���D�:�%%Q���8c�8�R�zݰ�Q�(>�s� �rM/�gx��:�j�Z�]�3@(ƥ� 湏�m^|Af ܇���H���dm��ݞ�:;~~������H�z��*�΀������_�r�.�|�!���@Qe^��-ڎ��؁}���){�˯��\zA��ь��F�����
g���p�
���:�Z�X*�����J��#@�C�E�|�7h�~���`�K�G��0�N��'���}�{�lv���P<���Z��zc>O�s6x��|H��k��62kw����R�]|�����-�t 1O1�Д'VH�7�+Me1�;8'M� ^Z*i�h���#hI�tC���F�ވ�����Ύ�,��*�*��C���w ��?��_(���J� �<j���/�F9v>���^�̫2�y�4�_��6w��Ϻ:؈���'��l��4��G�%y}�n:�М�!���f�9}�}�} 6}#��6�ڠg%�[J�i��k������m��>�P�yr&`C3p���pV)i���a}0�J��}��G׶V+� w�_%��^SPG���I�4��aV�I��UN���7��0�!�s���+>�Ւ����r�i��t�h-�U+U�(n��&{�UW�J��2���]�݄���p���۫���>��A ��j�](�������$�����I��]aמ��tI)j�;�o�2l�ਢ�s���K=1���sx.��=+�u���Xk.�/ʕĦ��A�<߾�бhWR� �S!X'F�Yw�+�ֲ�Z��r1�E�)g�`>�L�I0j��)Ҁ:�"��{P���8��a�9B��lujvr
�%9a.i�N��I;>�E�5��c��j����HUdP�T7L��n�q
C���|�)= �M���n�\Vy�RL�A�Ӌ����z��J���ѧ�~��]�v�o�˟^l��#sV%�`���k<&��{��MP1�|�
��J��A�l$8�t��r5����t�xo��F{��O��G��l���c�@��ԗi2���jL��QM���y�Y+W]uU/�?��)��d��mF�W1�
�� X�u�W��b`� b�}�.��Ҫ�Q�t���Z�10�1@|���X���5���)��p� 0�p��Q���������NBf�.��}�ԓRT��D�Und��>9U������9gO�UW�g'�"�[�N�����@�j���?ʋ�9~���S2δ_~����.j�LS&�����Z���m�4k�]w�]�ޫ���+��18��LF>}��k\0 
SsG�%�W�<��4�~R���p��L��t��ž��RQp-�
�J	g���>�ǹ���#��+������f1���Pi,�b���Wg ~���j��-�������㚨-H�9SUd՗�o�_��/��m"�`A����j׽�;����N�s'�����7�3 p��FE�� �H�{"��HH.6���£���T+�x��a�7虢��f��5���Vg�R�f��b���>g�ݶy�:Lj�,9)Jq�v"x+D�x}H���d� ���+12
ʐ���WN5��H��6����\e�P����7����S=MW����c�[�� (�c���L��>��z�Ii�=��tU�ŗR	3ދ��<���&�7�#�Xd7Mc1�>�&�K�i�Ҥݲ��ħ��� *��ih��{U�b�!|�ѡo�=[)�}�lwb�j@\��}��
�;1����f��)]�l�rukTE���h̋�[�ը>T)4�-~A�]T�Hă.��u,�[��:xCls�F��0;0���	�� �F�p>�y��=�*m�g�(S�F�(�OI}xG�r2����a�ޱ���y�,�U�6՘=���h�����vp�!�P�
�]�|ʞz�m���I�:c�&
�JqStPlT>e�j�A<x�	�VLH�td�6�YEi)���*�Arl��C���|���g��VZ���g�i�]w��>�b���	�\�ienm�{婴n�qz��Tд�-�I�trV��NO� f�X�A��?����TWk�[Z'��Ϝ��I��48P}�-6\��AyAh�9:��~�Q{�����.�����'�SOcF�Vc1�HFϵu�i�,%�zE={nj�Oe	��>���#�A��*����X,!�A�l���mƥ�5��۠�C�
�����}�o��O��B��n+��ö{����Q�s��:�vO.J��@q��cJR���{H���[#�9�^'�(��D�LAn�(���@�Z��G�)��8`�
����O8���1	��� mҶ�R��� ��N\��.�#���&��q"�X@[U2'>�
ߠz6SVA���$-���CZX���� [f*<�p,?\Ӓdb �Đu:�k[�ֽ�0je^�w^Z�I-*�$���b=�y�X��U��tu��OY'�5��)�2Р����uvyNЋ��|uoo������rG��V_<'����hյZ�w��B�~�Ⱦp,���#Mb�����$��?�+©�'j�zUF��;@z�6�YI��j\X�额q�Vۺ�b��ޚ�s��]v�U����p�R?�"	��Մ������5���$�� AN1j��O���H6]���Tii?a�DH��Zn~ ����V�(h�!XMt��z��v�^�<���޳c6�W_n��-�Ś�j���?|������ر� {)��HO���"�̠rV�5� ڢ����}�7h���T�%��`�mˌ����[n}~`[�a=um��67_�a�Ie&�#N��)=%�����n7�}J\�d�Mѷ����ٽ*B@*ψ�qN *�Yb�|�Ȩ5_���	���#E��:?D�{Pw��� �kt�?z ����s��f�!�e�v������	�N,�Ƈ&M���U��N�/<��\$�`%����ʡ�ngbX���Ǫ�N����x��2ܩ���U�^?��\��jh9��Y��^�u�l�F&�X�`��;��3�w�Xu#m����v�pÚ��=�$>�oV_��,P�aD�K�A��t˒֚����^Y�y5�O
�ϕ﫶g���ѫcAx���C��s�A�+���*�E]Bw�XuZ�Zu�lG9B�+� ����3�]&�U��a�p�jK�d�)�C���m�����+���w�����|�}�O�(�@���rf�����%t2B��B�op�0¦^-�:��I��l�\��˗_�o�*��Q��4��R��R�Y)h��~Jr%��,�۵!�o]�x�R�O${MT�q �g�}N����=ީ�NY���$���nB3˨ۺa�����R;���?����z�.��j۱����5�;rׯ�t��Y�~>a��A�+I���F�x_d����g�<�mO�XOb*{�D��I��ז���XPH�ة~��Y�/�?9xP�}U��X03�Ȫ�N�����rq���\�R7x_[��	臹wr��}�l�鿱���y���+���6=���漕p*��=�W)�}�y%( "@ݿݍ.p��K(�fc��}�y��(�m�O�4�7��Jm��/��;�����c~���,^��k�_c�-�1Cޤ�ڻ�~�ܯ˓�4�O},~�w�G6������W��N�ju"���G��fX�����o���g�]��b;��K��8����X��{���4�Q{b��=0|<��yU�O/�lW�>@��N�my#�h6�F��=7�XHe��j����@����6-�Vd�S�s�
x�,H���ي�-�O�V��(��|�-Λ�����|�^�����ZDZ-�]^��r5F�� ����Z������-�]�{F�|𵨓��pN��o)�Q *p%�����n���9C�4NF'��QB� ��Ԭ��KI|��+�&Jm�s��j�� ���u�sk��F�@x-�%L1=��LZ��i����'?g�~h���E��isI#\)e�M�D������ƶ��n�����o._�] -����yK6�`+�� ܩ�}l,�`)�����ʸP*���`�����a�^Oʥ��2p)�Z��T�c��I��`��*�D-�5�f��܍��\Wk-8�n���y{��OU�uߗ�|Ggx�2��D%0\ts��ߋ�e����w��'����ˌ��7�4�t�t����`��`F����n������Y#%]��t��z� ����D�2y���*�Ν�2����TT$�U+i]��˕ؿ$5K�6Ab�̅/�%����e17Mx���>�J;f���K�r�C�j�+&	ދ���jSM��_���H ��D���-u�z(��6��v��/�ZKlb�j;��bg��۪�vb�8��.8i�9cX�DuD7^�T=JK`��h�\o�r~��p%�㊟ך�{ݜcNY����a�e�Q�l��C��1�x�t	�xO7<��a :f܊�LO��rX#1�	�-*U"`x#w�_�gG���{��X�e�ڭ�u�i���b�F�Ϭ&Ղ|��LNs��KI#�r� g`!�TCT��ҝ���V���?ߊxLǈ������^W\qE�
#O��z�.D������ܞt�Өݍ�a�������'�r{r-�Y����2����Qi��C{������7��]x���X��C��7��K���:Ҥ�c&ʎ��wm� O�!��:��2����NR���.�kb�������� 5I����r��uXZ�b��ü$L�C�_��?�jfړ�FQ��=���_m��/9��^�Z�
�Нw�Ҿ��'챽Ǭޘ�fk޺j����Qc��h��<�Iֶa�z�O0XA`��H��0��
�k�'���A����7]�.�0Z���Du��k�F�J�lg�}v ��ǜ��*�' F%J��).�)L�)�C��Т�1��n��6�����x�w��gϞ���/y�/G�6�j�	��㜤� )Oe�~�m���.;�^��Kl��h�Fh��l��1=/a�|cґ�G����M���G�~Q�Nu��2����+����'+�(/n��A*3$�z�68鰓X���9ߓAx3Nt�3���#(�,
mPK,�6����a�fw����Z��d��"�i�����(id�ն=�ϱ_������7	��lۼ�fǏ�#��k+V�Xb�����P$�*�DMb��.�,F�RH��ɚ+}�c�@���7p
�����$ot��"���0�SS�5VGt:\� ��v�M7�ƞ�Gkr"(!��o*�;�������P5��ߒ�g��뮻b"旼�%��W�"ޗ�R�q��b��~�R��,�O����-��^�[��T���F�h|}9\r���,�c)Z���~�䋤c�b�l���A�������-����v*���>��������Wx]�w���뢟n�����̆y��,� i��(z_�( 0^bj�wۻ�h�O�$'��1�O�Լ��� 9���P¨T�F�w��ٳ9zE|��='���/'�ru��@Y	x�/8B�0$v��/}�KG��e[�� ����_p˔bS Z�ت��涬`��q�0����m�{�����}�=��S���J�̐��ΰ�$աc�(�Q?N:��P���J"�s�=�^���/�rs��2���>�у<!�d{����)�ͻ�~9�V��f�R�ӴV˔�?|�)+_W��Zf��"~�x<0D���6�1/E7mǪ%���K�r_�Iu~�si�K���dƻ~�`�+�8�����t`��~��n��Г$���uJ��-ñ<��#�L���g�G�17�s�OJH����~T�W9��4b��Rq�T׷�h��G��"}2��)�I�[���Cf׬�J�����w�"�|�gon$݁y���3,1l?��'��R`&Y&#��V'�jWVs���;��*a,��G����0�m'����l�D˶��;������<RD+���^�M��z�z�9\)�õ�R79��L���J]�q�6)@ə��ԗ#:�{�qn��U�P�8f՞��X�����ʓW���fl���:��`ɔ[���a{�5W�A ��x��hx��I@'}.`�\��܋_��8����IKW��?�S?��cء0 ���cy0��a�<��|�3C�/�wa�,����w�=����c&����2���aB#� ���{�>a����G~z|�R���Y��1��8�(P��n4��� �Q�
��`���{@8U��r�23���/��[� u��Ja2�ݜ�qaR3�}�n��e�}!��ϯ:�=h�ő�d����'$��t�'���Y�U	�>�po��N}���ə��ONTs	�q�����Tع$*�$jb���[:�|�[��{�id��)�r��$΅X��m}?��	�pȾ���>���h8����;ڶ�:�\{�tû/)=+ 2�06���	�.��(�mw�����k��Q5F�+��2�� 0�l���1Q���Nػ�o���3��y�e[o�˽��^���[qΈ����ΞC�Mn��WLȭ����~$}�~�;*�����q�u���9�~~:�Evm�nZ���ޭ��׉zǩ��x�7�Y��?�A/���׽n�v�����K�
?�^�8�Z`ﭷ�:탹9o`��cp>�{ؐ���
7�|s��*8�O,{�XjG���� ��r3Pzn�|�}~CJ����w\|�nL,�������7�G�%��q�q���"`�2ep���g�Y3��!�9��J��o���1	=����~f��M2WT���J��q6<p�C鯾�t���:�6v�����P��l.�n�A7�[k)[�[7QF���8�=]�p����h����r��zʠUp߭\���y�G��zg��b
S{l:�L��섃�g&���ի��,�O�1}��ۋ�@����u�r��9��m����"5�0;n�`�m��n��c���aTY�)}���D��kw�-����&[l� ����T��׋ 9�4�7��w��&���5��0 �[o��m�\��6�ݥtp�ĵ(ӃS���F7=`����ݕ�3wB���X�N�d�J��Zݏ�M�� 7`����������;�i�F�"�Hl���z9,���T.	��>���旁p �9&����Q�;�nq������4����@t�w��/D�$�(�iYII}f��er^���"]e��`~PU1���y����|B�LRC�h���kl�	'�
d�,�
0�c�-�&���Ғ;HKt����u����v������ݻ���t�=/^9�m�	g�h2]ty�����t�iAZL"o������̛�*W `��g^��l�) w7gyj�/�NR�*�<��@��P��T��!3D~�F�ϚBv`j�޺�1Q1P5P%>�&Xiky��"==VǚŊ�?��פ)2���e.�.=
gBh��X�2UҔkPڽ�NS�?�$?+�^DƵ�z�����u]Ϝ���@|� �VZ��=�I��2�k{i�����d�ʢ��]ߠEX�]#:�׌���*��\r��bV�̒`Ɵ�ɟx9X
����o�?��OA���� ��� 6�͑Z���'hͩ�3�������F{��Z�n+��S�+ƝZ��ˢ1�㼳�q���4D�q���(�VC����x�)�iB�c���(�x�����L�W\�R��ot�,���<Nn�Ml͠����F�&Mz.n��0�|v:�HJ����:�w�r1�k:"D���@7;���C���ܸ����x4q�Y6_g~e�L-:)�a�c�Y��ô�������eS��T�t��j�8�ndǇ��d�� �=��)𬨦P�h�v0��ݛ��o��t���7�������0�qݜ�6\E����X5N����6�������^mV���TL�S�M@�aX�g��J����4��4[+#��Cs)R�eb�k�ήk�B�6�� �:�u���O�{��g�p��X�Re�0F�$��5�\N6kM�r!{ՅM�?���1C�5���x�);��x;e�h�9.���bn�k��֣�!O{2r5~R��f�T�Kf�h놌�C"�����%X�i�$7�$e���&`��,��g0�^{�4u	6~C�����+L�`��` �t��m�:��al��Z�r2��Fo��G�������j5L@�$���ÃE��]�yԱ)p�=��WC�ѝO']Q�0�����`g`�"?`�f�[wh�_۠��R�/��Yh��d7�7��)��� �ڌW�U�&<aM7%(ޘl�&-���U����	�%�w��`Ǌ/f*W�'��@a@�!��+;(�
�^#cR��D`'�\���y��I�Z��ʺI~�2���r!����*���SG�y(_1��?�����o��-�T����y�SGdfХg+r�9('��9󩗳#�	sϵ,-7�l�����^�� �XTה�C��`q� l�L8_C��,�&�ՙe�u%h`e��05��Ɠ\�&����q����&���Ν�Ƭ7�wҀb�_z�F���(�!�Yk���E��/�y ��d:�S��׌�,�M߃�|/U1�ħB��^��ċ�T�Mv1���������X@@��x�K_�{���Nf�	��Wjة{��>jU�~�4 ����f]�E$\�i aDv3d&��sB�$�`�Y1/GuB7���L�z��1-�E6>�'��I��?���/��/�Q�����漊���G���ƄMjV�M��M=F�0v�YXX�L96X���&u�Ė��s�i�S���ߑ	ov�0��]��ls�曞좲�Q��zn�Rf���-:�ڰ�ONIU"���F��0j;��Rׁӯ�0iR�9�7V�:C7�R�Ә�w�^70�pV�{9��N�(;�r��4�����{���^���:�(�iH�s�� U�
�E��`�M� �|Î����V��ͅ�7i"�f4�;�j`�,�,g���,��<S��l[,-�=@��ݘ�h��g7v���|e��'��j��>&����h�NV4�ko��38�βobc.��q���zӨrF\����`ves_u����m�ct��p�MZ�K�A,?E���ϵ%4�����k���{DǍf�F���w���h��3s�����?O�*C�t< �m�N�U}+c1���fl\NS��q�{] \�#��S�z���*[Tl2r���r!Q:�dZPؚ�KD�����U���~�{�s	H��7���Ƙ%86 ���񌎘�9b�p��G;��!���3;�\-��C��iV�`V�=�W�t�y��w�!�`b��k�R���s�Ygo�EY90M�{Ӿ��^�*7�tӷ���t� �y�c.H^t��ڄ����ܕ����w�K�R�������=�
��t�y;�y{v�]����8�ԛB�`�n�)�{�����t`ߡ����vl�k��Ҏ��}�:3��B,AG��rz�����ޞ��=�q��V��9��L�^r���p&�H�)��BsF=���Vc!{�:�9;ܹc)]u�S��h��Y�ày���r����ӏn����ђz��+.K�G��j�QҘ�"�{�k�������<����5��\�']r�cz���MtG�M���O����v�����a����.��ϑ���ݬQT1���V�������}����;۷��'^�ce��j�*�ܾ3�|]�s����[��H�:5D��ID�����[�n�N�',gg�g����{����$&�:�C�ػ19ֳ}�N�\��I���1I���Xh��������+.�Z8#ӧ�a���}z]�|�h~�[�?�=��v�m�m�3vs�� ���MjB���AP�� e��Q^���s�Hm�B�򖷤?��?���w��镯|�w��H͓�Dq��(��у��o���FI��ǋa�J�[����E�xvO3��qV�j�*5�$�9��$�5���`���7�"=�9?al���*ؿ��vdlhh�뎝+&��������?�A��m ��=�)����
�L'��Pڶ��:u�E��qR�x)������ޟ����r�������}B���~K:��mv�5��^�Nfs�%����t�?H��;�o*Lc0�u������ғ�|L�/vlْZ��Y+OVӶ���߹#����?��H�{�X��_v}z�k^h�q6�:���n������O����L+X�k��	�����v�*���t�u'��c�q��*>�_|��?���j ` 5�ϯ�ӿ���O?��K��u _���<��csxם��o���j��v�];�W^����/{zZږu�uX�v�D
��߳绔�������7��Z����7���ڕk(8�� [[?���qpUv��y�_���]���²}!����o���9m`�5[��m��5���(�/~�o����-�y�^�����;�fK�s��.t���瞫R��ۇ�_���TW��yn�L�7M�ұ�l�i����d���կv'k�+�FK�L2�@9�d*Qx-B�ގmM5f�Js��������@�@ �����).�S��uf����ɍ���t���Ä�Fe�0Ĉ���E�A��ʰ��7�t�O2C:���⃉Ԑ�W,;���#�!�����[3�ܮ���{�8�y�##g(~�c� =�����Y����t衽�k����M���1�]|ۙ��:Bǘ��`�}֊��e��iea�30:�P8{q�L�V�껲��+7���g��{��ťIZƙ1�a��@���R/8xwN��Xp�_Z�Z�6>ҋ.ܕο`[Z\�}���gυi߾�n/�+�}�bڿo�m�����$j瞳�X�Yimx���L�+;L���}G�l���x����s�MȏL�䒦��/�s�X����<ώ�fﭥm��2�ٰcV�%w^��s_ ֖��=�3��ڈE�w�z:��rmt8u!�Hq�&�� �m5���`Q������Ε�K�;w���&������G�`���ׇ������w��cǢ�k*����{�=���\��=hb���d��c�K�&8V�wl%؏����w���0mhl���Ǚ��si)�d��k"��57'�Μ���2G;�1k���dSM֎"	�j���s?�s����8_�?��F)��Ϊh
%y�E|_Z��R�-X@M�2g�8��j���h���wZ>�i�Eg\�L���.��0�
fw�u�1��א��pF� ��rSq(>��F��D��]�z�� ,Db�9���w��_��4K2غ\�X�Ԑ�@b�ǉ]G�F,p^ٱ����4X\p���]{�=�ܛ���Ϧ���<|�IO~\��T�ڝBkn/���7�wpݓN0#,���T��|�[���HKۗ�EoOW^uYڱۘ�;kvHM`;]��J���T`|�onM?�����祧=�t��%�\�9Č���QV�D�����Ӿ���}S��������fl�{nK���µ~���� V���i���ih�S7|5�r��5�S��.�e�ԫ�'nӦL"���@�+t0؞�����w��}[/���������v}�=�^�Z��YY�vC��m-���;�}�>����uO�:]xɹn*@��:i?�����:;�*ZZ���7nN��v�k?qՅ�k���pSHi��2��",Uǳ���Nnڿ�7�J7~�oS׮钋/HW_uiZ��w|���&� 4�b���?���a�f�������A��>��?�t�y;�ֽ��y��Y��<T�eS��L�uwJrM'[�d�!b�)l0�}���;  �$e���ou�x�^g��������<զ�m}�(㖡��vk�I@Dx�v��=F�7�҉�[���舜*�Y2���w�c�w�d�r�25p�y�v7C�(���Ka��FdV�YV�����X�DH�Ƭ�A�N>yI���P���*��"�b�����,�}`�1�>ے�*<����=���ƺ�����ϸ:������{�Ys�0@XXr��`���rE9�y(�G>�����t�w�sU��O>+������W�pj�d�f堟��J������o�f���{[��M?0��۞^������Zc���3]J�Rv9��D�Ů}�a��?�����|��I�Ȼ�yOO��S�s�n�Kf�\�R8��������������L�?K�ݷ��ql |iz�~%��ϼ8��Y�z��׺�I�(�L�կ}#������������Q���_���o��0�N��~�f��xT6!][/��[��O�����X&�~�^�^��Wÿ �&�lnM�3�<"���q�������|6����M{|�M�}���[��7�s�s�	%;s7��ܷaZ
� t!撾��/���_ߖ�}��3YL�9'���_�~��ޅö�g�~���X�6[�ϭ�ݟ��~{�䧿��eb�����_}ëҥ�{�=��L��n�� ��l�;�\��/��j�F'?"���l�z�����Nn�U�H�����D!m�������l6�p��}9�-�Z��3p~�*�5Z>���mm�}�<L)�j�i/~�En(?� 3����R�)+�4�a\��&��ᆙA�Y��|�C4�¼�ı�I!�ɟ��������n��
2��Um ܊��9Fu�̈��m�,���ݾ���s�1��N�}������ie��tۭ&�׾��t������jKS;��Fͥ� 	�1����}���M������|���L�_��t���9�r��]��.�[�X�>��/�>�۟Ɗ�b���}0H�x��M|��Ya��	�*nO�z�uS���nL��vȄÂ-�s��>����g~#��k^a,|��q�s��hB=�ή��o�bZ��������a��ᓷ�]g>]���`.9�Ф*ܴ��Z#������_�n�X[pG�n9����䟦�_v�;��3��L@.��u�'>���?�t�@�7X�̯?~���%�=1����gɜ��s�Y93�&ﬤ[~x_z�{?����E깣���t_z��h���ڼo�=A'��,8�h�Z@��u2}�+w��i}������K�Y�??�쬍���������7��`��JkƦo��W�ܟqM-�h�?��Ϥk�{F��1O�}�͝��f���3�:�&,��)�O;A�v^�5��[���o@�=+|��/ RMt��p�?��ϟ1�g	^Q���"ܐ}YF� �F ���O�[��F���َ2L�K+���w=���ȷ���/В�M6��cp3$[���H3=I$�M06�����G?�Q�j 3�;��_�r��}=	�@�H��I�A2VU:�!��Vs�=x�����T�r�	�����z�(zg�mw����~�Ύt�}�|���~�m�o{� x�c�z`-=��aS��H/~ɥ�{\�����c܇:���0=�qW��.�A:��!b����t�}�l��I/�k���.cav��('X�]w�7 YN�\�Tcaw{����ko��>��]隧</]{��y��84��P�m���xMZ?|K"�r��NS�/J���~��������[��_���-=���٦��KLwl����-y�k��ք�!�0پ�"�d�Ԙ�iI��, �k5�}h���K��ړ�x��{�y_|�9i��a�׮����_n >rf� ߷apv�ѭl�[ץ[{w�ZX^��`���M�S�v}z��c���y�����G0ƾ�.{���os{��2]asp�	�U�OI/{�N[{�j݄����Qz�������Y��'<)=��m���*�g":���g���j,���RK���w��Ɩ�t��ķoK�{����9w̕M���m��~� |��!�2f�i�9
ႍ����'?ُ�}^����U8+�Dż���o|cZF��������	����:�`��{�= ��`m���D���iˍ3�'C���R�}�.�8�\�X�*֝7���	��H,J�1�0gl=H���8���JkH4��g�� ˎ�0�hw�)C������8�$r� �
MS�����y�����_�m�/��I�7�*o��u����)�f���$�c�Է{^Z�Ą!y�}gүy�y$l��6�!�xki۲���*=���LO���.��xW(����ܟ|I�'/4�u���.�n0�=���%D����e\�F��^}�3|V�����H{ο��m�1�����Cv���HYIW_�ܴ���;�{�%��/6�Z�ݻ.N�{�����Ҡ;p��ֆ��+�N������v��f��"c�}�����r��@���u����⍴z���򫍑ߞ��w?�g���>���i���t����=+�֧�&d�<P���g�8�oH��zz�ŏI������� ���_~��ߡtnS%�X`>���Dx哯J���-����<-\c������'�N��T^�P�8/p�l�����g��o��w.���g��;�\uͳ��������6pX.�����级>���_�YyT~k������0ը!�0�#��+��}�2(����I�H@�d��s��9��h8�L����a:w��UD��}���������@(F<�D �+;��g=��6���"8
E�5n��g�
&�����d���.��ff�X�Wǅ�������v4sB�l� ԱNv�J̋��^�Nھ��OT�"Z�ӵ�ޖ.X����O	F�I�=�H�];�2}�C�P/K�lm{eg��Q{M������3U߫XFUM���6u�0-�c4,�Jc�;���o�(������ٿ9*킁ނ�gl�ۖWҶ�(���z��⒛P�Fa�E?���"a�Z�<-~y����bJj�d�K��F���a���:��AG�3�����+9�7�ذhs3�cO�q�� �ޘ��E�@t�r���X �Ѹ�����\n;ǎS�5M��������ߎthx��υ�<#*k�vb&|�&��\^X���HR��wβ���!*�fI��{6�6�E�ڗ0u��z���p��g7��j��/,�i��0H����ǀ��	��D0c���i2J���f�q4�'�/�Kc>�7��f�JS�lDՍPsU8GЖ!��髮��q�^B@ ,�p����O|�΂�5!x����c(�3�p�IB�.�c�2�����B�I�P�Vu���#sC�����%7Ex"Bc��#
�5����F�t����sD�{, �� �08�U�v�D�t��*�]�G���މ{��ȹDכ'�g	g�VX��.j2��6q�==��3���Ң����7�j�Q�x�3�6F��p��M���9
Ï��f����
����g7L�+��լ�z�_� �v[��67y�02b>�3#�k�G�NuN
���^���4-�H*�q�l�.�q
/5J�� �g�"�n3'-P��.���Ǿi�e��+@{�5<:��ϻ?O�i4��s!�_\1�p���� >���Z��3�e9���mv���|�x�:������{L{vc��2���Mx�z^��0�%7I!	��� Б�6XH�W�=�sm�p.�^�Jj*�?���I�	oZ�[�#�b�c|��͆$ŐW�m,5b�#���/8�&�S*�G�:Ų��=G�l�_��צ�'D4Ci�¾W���FŨ;���7�JE�}��^��-��0 S���L7�B�Q��6�P&��u2g(��RL^&�'5G��r̓���[�f���L��@Ք�TA�"���ey��\^s��Y=���&��7��sX�d%Ϥ#���d�qΞ�S�F�I��$�.�!y߰�S{!�ը{���+]]��R���L���U��笻^g��j.%9H
��f�E!��Ef�9�?98�zJcAU.��Q����]6��P�zmfϹ�p��� �N��M"Y��P�&��g�7g��q�\gѴ|ϥ�X��x\n���{��)�#B�:O�����:.ܜ$�Ru<>2���g�t-)F>�0��W�x�)��r[�[zd�t�"G1�U�u!��a�؇a��F��D\�Xs<H���`�0f�UL{�uaNf+B�8畣�M�n��N�iʏ��V��*�b��t�wѝM��8�m������K�P҇$#�JI�h�9�!G�	ozϙU�+���:);_:��C���R��%|�k=�^���T��=���uP$�"��!�Cf쀵�NYR����E�i鵅�^��KF&����L�t[��s���n��5*���-s�aS��;]Pns�j���)�$|�^B�r�aO�����'XpG�g5� *z���{�lm��IE�β� � �e:����R2�:ɵu.���z.VD&X��5�&�'�v���GUj�=��hrHk	{<�Wk�i��n^�Qo�4ʢj�q!�M�CNZ��Ir%�f.��I���M��>��p����h �n�
@-׻��0�#{�.4";�N�oI	�x�D�M �֬���1q�""���QvGͽ��l�)����"H.�2�4dL�$��r@�ט�[��0!;���R�o��T����#���2���C3`i")S�i���)��M�t��u״�:����sű�5�Nw��~Y�e"�k��s<qSϠ <+�i&��穩C��y�������۰�:; �IngT�3����=���f]%r�G_c^S�x��47��*�����,CBB��r��=sM.�����(�.��Y�tfdE��6�Ԕ���$�Y�^�jf��M)�
g�.�oM� �� ��2w���E:�Ng<7��2�\���	����!�^
�!^��>�4��dVߝڀg�Xv�G6#��lLcDS�!���Mْ1+f�>1<3D�S��Ĭ������r��*�̖9{M�mU���@���p�Fs��#�jK�n�@�����~�dU����=C�EaX����j��+�h�6��eS7b�����N&7��VPPʑ�C�̒�q�4Rĕ���}�r��\X��ISƱce����*���2�z�9/�6<��Cv�?�l�g��F'��>�s
��$�G6���#�g@S!rŃS��Ռu��V^�`2]�̛�O�z'g���Q�l�.<����KN�0��"C���^��9Fn2��{^�$g��ba*�>q��J�Q�g~�n�/ZC���$W�΍�C�GwT5�N=[*����ts͸)�T:㧤e��k�*MKw֏l fDBv$��~-�[<�2��%���������C;�k�i����`g^�ٍ����p���^������n�*�#�{a�5)LD�� ��0"�̈봰H��<�=/�΂�$�aE���q�e��Ȍԝ��ȩҶ���=Kk
�tHn�$�  ��v�\wOz�o�d�����>Eo���X�d X��r���r�m�y��>F��g�ts��<8IdP���۵�^�-<��	�����٨���B���Y8"ȸ�ŉxo@��Q1�M��XgR��}�����$C���:^"?���gsI؞/{?ޤv��3|�˜�[,�B/���M" �t���\��>��T��Ft����\E��M���~t�ML���7lf�tt�y�8�7�m!u˦��x�S���\5fi.��1�{HGf4�0�]Y	�cz	��n��9���.�Hɶ��7�@PW5�u��,m����VC�y��C�4�����HGd��>��[o�^���ﲍ��,�w��^�|��hG�1P�g2^M��Fڷ�J_��_��ݹ�q��gv�u��-`�ݎW�"��`�5c���ލ�o����`��)wi��<�t[���Kw�������������/~m�T3�k=s֥��͂&r&���<c�;߾՘���!egdٰ�ƖI���r�GUӕ�������r��D�2i &g�i?t���3�MXw�q[��WK����gբ��ah܃W�릛o�݅٨��B�*W�-9h���D7�l��6ގG������ʴ����}�f/���V΀�ٴ��g�
�1�Y(r'�J� ��fW�ą%C��n$�C�	9��7�!{w򵔷�#���i����XA�N,�m$w�͔>�ZβK�o��7�?�#��B���'�Kr��S�1���Q�ěUL��l�
Q򇘵� ��$][m���ǅ���ŏ ����r�ވӀb89�=��m'X��7��8�}��Й���O��~�L�W�{熬�e�z8ruvu�PZ\�xA����� ��>�ZԒ@ƌ�{�e���}���l﷍��[nI��r[�� �9�P�N�A�����%�O}�=�>���h.�C�����Pbp����v[q�{�M\{�A���#/0��b�������?8:��uS@��e1[�5A)OB�;��d��羐r����jb2�%�=�Ո}#E��[�F�~:D��M&W�9S��Yh@���w�|��/ _�2@q}�o6{��>�;���Ye۶�Ё���jj�i�K�n��{䐔�FԬ�X����~��x4I��X�!�N�\k�Z0��=':�):b
��4j"8����S��^��ь��{1�WJ�!67Ɯ1�Gژk��K/;Xxo�D0�^�4VQ�;jZ�$w�岀S�sa�!`�c�SjL=>?���z�hS����rn��x8A�ڜ�&9�id:j%M�a�;H����ZK��VL|�uK[���?�O��G���x�[p7�GM���a�p����Mf��z����7V��q5�~{#��z��Ta��\��0�I!_ل�\���jԉ>��oz��٫aj�7n|�e��a��ٳk�Xp)��3ہ�����/ki�ӧ��X��ςU�@pv����LaD���h�Կ������Y��r���5N=�ǽp����QB�"F�Q�{��*���%�b��5?�X��GS��Gp���'�0��������S鞋w���n��l<R`���Ю�|,�,���@�Ld����n���s���]��Un�w{����Z����XSfԜ{��G��4��(����^���Rs������h�ߏ��9 �@�q* �l��XI�A3��b�0#2�v/��1d��w:!�9�ܖ�N���o���jb�Vj�!� �~�匓ж	=���ϑ�2���8���{G����1�9Nd."��w���8��j�ۼ��s,sq,�u�A�I���h�TY\�@Q8 Sf�F�L����`rصK���6��T���U\x���G�>ua�p1�!J�^�7-ƳՐ���+��x���H�=/��h�?@i3�c1�̘��N���@|+A���JA�vm5�5/a8���hю��=H���1Y9��J���#�K�e*���Y��t�h[f�֖)�ũg�ոWl�
~��s,6�;��a J�8�iB�_�x�hr�iYu��;N�p9����X�D۩�՘r��9��\�����^[�c Ȫ'#�nd�1J�CɄ�* �9r�+�͜S��G�r�a߫�x��	�ˍR�Dݔs/s<�іMц�Ր݇�(%P��TH��yl��؝�8&}��'B�[s�Bu2��p����6��.&+��-bHk�DA\����?"w��[�s�#5��L���#���b{��%_�t���qH��a7V#Ou I@��,�*�VC�+7�\}�Y"� ?��0�}���ĉ>��}��sr2��h]��:����k`���53d���8� �*��QR��:7"u�Ȉ	�Ĕ�b�\O����֖ �+=Uc�
h�#s� .%*/��R�LD^��ƹ)�@P[��XR����%k0a��8�{3q���S\��=q�m�':��$p:��cqXI;;U�hL�s��#��4 F5���0���:�I���d�M���#hSϜN:&����$�P5��Ԙ�����ܔ�Ʃ�	�`�����M��L��27(^s�5^(l�$M��q
 �&P6���ƞ
FTV�TS�8U=����z�k_�R��`��_��t����!�>��O�}�C.T��q*�t�c�j�=����od���Þ<�3?n���xQ"�e/{�W;c��Έ���/y�Ko�7g��Q  �B�/������Ee*�v�, ��(�IsO���/SEÈi�q��#�aI���^L��q�k�����E��7��b�X$�@8&PPY�E?�'=�I��Y���4I<�K�xz�=�)OI��|��ԧ���˿�I���y�s�?���(����ʝg�?��������I�u��W��������I�f����1\MQ|����E^C�أ��1������{ ��C.U�2��DK%lm�0ܡ�XJӛ��*��6��=��t�嗻$�,@�_7�D ����(ō�l���`�0�TJ����C����5,�g�a�L�����O'Oi�qB\ęqf<�" b 2&��U�J?��?�c�d ��i��	�!���gz�`uw��{���2Eo�c�; ��=�y��7���M�Ɯ�p=�6�d�N��Ki�6r�
�4h�y������IP�O~�4I#$��!�)� 3�8^��:8c'�6��1 �4}�+^�7�g~�~�M0pu�PP����A~$�93Ό3����){F��`��׿�����>;;�tXva��x!}��캊C��<���y���M|Qh���&�NEQ����sc��pq�wp�FnRࢸH
�sQ2l���xj-��M�LmF���,���V:k��1; �L2��x�~�����Z�r
%�q];3ΌG�P�����}�5�y�)Z1L�����܄�S?�S���!E:�)8��� ,��"*"Q��`�;ǀ$�XD�:��&d�����jR���b� ���L>mo��I� �0]�$�I���x!9��w�N�����i����X�Vc����[aqL.��n�gƙqf<r��%�e	^��pѾ�����zM]�g��$h��`V��g��2-D;/�rNp �[<�A$C�6���	�I]vJc����;��p�!@G�MIރ�"q���'�C *�	R�/�5;1��b���Yc�A�5����s1�?�3?�Cy@�p�p���g�?�X��1[b����L� ����ڵ�?��\	�k2=/yP��l�;�+0G�#ӄZ����t�UQ�+־�&|ʣ#�bSQ#<��[��x�ށ�2�L�)�q�|N���XP�C�d 1�)�c�m�&��_��_w�x��L�G�>��Ϲq�@��Q���V�*p�錝��83�e�h���a����T �������{y���/Т�  ���A�wԵG�l;H��bBS�#�$��WҴ����pܩ��Y�+:N߉��瞻��7����2R���
n�5���q��7ߗTSz"����;���xA�U�.�G)6�����ԣ�<?���)�i�S7�+UD0w������^o�Xo��\������vѣS�-�H}����K�������F_)X@��W���t�7LqQ�E�ٖE ��M�7'ƫ�f�2�x�F���ٻ�'��EK9�q���1�=N���M������~ћ�E��g���ȉ�Y��thW*��A�}��w)DV�7��Mnfrc�e�Ek��g�ԤF�^�;,��i���k��m~;7y̽��鎿_W['S��c>3N瘷�Ol=�e���"K�c�����.7E��oH/zы�������o�qjj�o� ���
]��H�x�j�����6��P��贿�o
�We�Z��Z.�~�u8��skn=T�Ͽ�)-W\�nP��$V�<C��&A��߀,L��~���CJx
���u�sI��3�ڞ��8��3�f#��4�̩�*��i`��������W�ES�*��)�K#�3��8]c��?�<�Io^�d��u��-N���L�����b��a�Ҷcy�؊(�=��4�A��{D"����r�m���-A�c��锹=w���`��x����=�t1\�b�f�����\��4�T�"1d�����=�d��yX8������Όy8��:����y�{�u[�W��zsQ�<�Pc� l�R4t'):�ku�83ΌS?�懶Y�h�y�8��&<�'��w�=&HH�˷���C/x���2?���W����>�'"	��>�a%��=*��\:S>�U�F�_������M)D�-���\��rp2�K5�Q�1s'���*{EG���������&�8��b�����.[N�Zʠ�j��g�
UΤe�\C��(+��f���j��jG��3�Q��B�c^g�����>�>�6T��?��� F�c�P�� :
��_��+���%��MR��b�ص�+p@X�h%��!�Z��g��oxksĠղ]��<eY�]g�L��AZ_��[5�i�t��p�ܐ��	l�HX.�p�v�vM6c�$��%6�	X�R�e� ~,C�Y��1mne2����g�6oB�wJ�0p��:�������b��c>3N߈���f�Gc�G�����T�:`�����w;�3���%4b0 ����5`�� ��Z��`�2/0�a��e9�%�q8.x�5t�3֝����~ԅ^W�l�U+sm`l0O�}uX��^��Û X_Ib�
��
�}�P$1w�,��!;���m�]~�b�T�GP-�m��)��+J�#�i#cq��"K�c����ek
�9�Òs7\�Mg��,���3��3�4��bs�&z4s��z@�}1ѱu*2WE�0;���o87��%��5@�$0�2X~���*���1Ҧ{�]������5d�I�i�\vG��	
�$1��(���?HW����(�zh�n*'^ �j����3��"@��"�H��*!S7H�5�Zbk@� l*+���/v�ü<�R%�;�1uʀ	* �1l&a�*���
o/�tS�-���t3�ٙ��1m�әqf��!�Nb�G�cq�EU^�SU>��p���'{���wyf�.˱j�@Kam�0��`�I�>Eq� ��5���\��s�po��焩�Qi	�rFk`C���|��_N?��t��d�ét��3��S 5�����_���}2e_Aa��+8�G>��h�X 7�:��ɐab��'��>�չ��&[f�t8�,�ic�PZ^��h������x#M0����,E�Y�1����pL��N�tf=��������P�6������S9A��=����L���L�G֦��0�ΜxM��暡g��Bճ[���u*���%�ߏ�i9�֔3&��S�RϺ(6T�QlI����[�T����Q���\߉eY�7y���b�����o�yf�V�<[�}F߈�I���h>�-.��0�;Q]��6�G��BW�����ǵ4o}i�D���*���x���Ҍ��Km�M���	u�͂1� �	+�-�װMS2�h�M�>���2u�NVۛd�`����>������!҉UGX7�E�bPzng���~��n<���zP*���u&���"Rڳ��c�����`�t�[V�k���0{�ũ�����d���R��U����Pw=�Mҳ���	���`9��Ua�f�<|(�y��k4W��m�3��D��6��ɟSP3��kk.cXN;����q��0DE��,"���Q��q�ц(A�s��qbcƨZ�dc�dLT�E0�wb�,�������lϟ%�d��rZ�
i����k$�g?����磹��IQ����9"��ׁ����j�;�u��p���k�5'���	J� S�G���I怈����b06���ߔH�%0)��������	�;h�C��N�8j�e�=U9�����v�^z�S�꓃���r�jE�`q21 0��=��J�j)�Z�)<�X0�I��j������l�?h$�(��I����sv�z����0���4Y7 6��v�^Y��tO�p�KȞ��~z��Ҏ�.rޘ��λ�I��E1sv(�$n�MϠ%��_�U�aH����<��z��Њ��^��o�TF[[Խ�Z�uEO��'Q�n3�M�v[=k�|E�C�MM܌�P�5��ⳬS�[���j�<T�J�V��GdB����D ��� MZQC�@=G�T��U�a�1�I�K�����c$�T�ڶ����h�k�<\l�B>J�ҵpm@59�t�|����<��`Eh@U
S�	������o��?7�#!%�*�V:�q�*j�lc�䅼h�nf�D(�ݻ�A�e)y�Z`L��j ��&H\n��b�I=5ew2e�d��L����������mS�a:�3\�����0m�Hc�i�L�o�;�L��1?$n����z]S��:�ԫ�>�*�Yl��`p=<lm渨�����.��{b~����o/J�#1a͹j��D�>��f��jck��Y�X�|Qx�"Lb�z�\" k=H��њP�n	3�(x,�{�f���	7�Pe�X�@�)Е��c��L	F��ya��9��F�>/� �}VM4|F�s]7�M;ZC�5�sH�E!x2� [�Yb�c߸H�tj��� �-�^aN�_�������7��y�w�|E�TSq��xtsD�)�d�OV��^���Ƃ*�M�t��܄<7s0^-ˈ�$Q�e0	T�GRi��q�yO���g4.�gK��b4d��c2flG6�P0 .�1f�I��ii��a|Ua��h@�En���Y/���{�nV^�s��$�z���,7f������ʓ��`>����N�P��h��L `��uIeBj��GtrD6�g��1�R#�H�&�X5jM�髽�/�f��\Q;�J�om.]s�=��hֶ�1�:�3����Q����ɼ!����(��֠��.^׫=5�v�A\x"㎎>�qt �[_�2��������K�A�F��/ӵ�=�t :�	�C#�<�u�s��^�k��jFDavl�i�>�z�2ؕȎ�v3��Q7��Ҡ���=(?�
*��D��ő��a��E�h3YZ�L���5ǖ=O\�Q��h#/��*��Be�W�lA�vX�^����~�<�*���ʩ�%��Pc-��0e�,<dc��R[���b޸g1Xݣ�����Rs��m����ܺOƑؖ����D{�
�G0��#��Jz֑-���)@����5�_	(��~�di[0�L#�D�b�1����������"���~#co3F���Z,�=�q^%����H�p$տ�^۔��q�g�&2Ui���ccp�cQ9Q�eQ��פg�\D|���N W@�-�����x��=#	�h�kk���p��V��B7,<�A����ͤ?L�����T�B):,Z���iqkB��8��c�6H���&XFcy9gj�_~�1��������
�#T��Sy���T�̀Aẜ4N��ɣ& ��Ttlsv���y�����]6�v�T/چ���0�5�V���5�,@�T��E+�)՜��(�E��&&�+۶Y4*m��Y��)���H�"�^ڂ�k�����F�?F�(
�m�՚��x���<en�YM�X�����^P	 1j�p�f���5q�<j\�b��]ku=Q(�AYj{M귀���6ؗ1��D�� k�k�ه��_p��ڋ���Ks�&��7�)��s��k���#�(��υ=*&K��f��ؽ��Ә@;lʙ�%�WLL�Ɇ���ʪ���V�d��MK����~�Y2����<�ԫ|;e��~�I �669���ML0�k�m \t��r��oRx�v~�H�$J���.a�ndw�m����[�M���juu�Ȝ��	���?7=���{|��Ճ�7�;���cr^g_��������~&��{ -�=%c2��l��;�W�������=�g"n�8X�lr���[F�%������g?�m�b�Qk��]���Cj��72�ig�V%�Mt�I�s<� q�j�6B��vZ�A�^���CmU��(��@0���2ma�� ��ԧ|>�k��>6!ҷ�76�z�����tŕO�s��.�����'n�tZ�=�|b� 	��]=��\͢\d���(������F�C��랢�"ڡ�}��s\=��@����A�	��)tO�c��?�HĮ8�G[3�aװ �ș�b6k!4�����4��u��ۖ����I������P��a�9�f���΄�Xۢȅv�����\����l��.80�;������NDWTv9��1ݾ���$8��a��G}5�cM܎'n�÷[�O�:A�c�#ۈk�i�9{Үm;�D޾���Y��i8)����7��ඥt�TK��L�F��P��?�d;��h5�}�Y�
WRJ��mz���"� O�Es�g)W}c���L/����F5��c#��~��
9��%��h�I��1�F�$��E���(� ��Ħ�&�/ ����v��J`�	׳��3�]�3'%�������{}c--��H;�9�C&K"q��c��ʆ��8d�dt�������	���}��~>Cy[�k.�i�N���=�ԥ=�~�N-�����5F�������8M5}Đh�o�i��{m�,~�mW�Y2~&���L<'2�nY�ug�Ņ�-�������w��BtDck�EWgV�����N���q��#n�u$����M�	�i�$8֘�0`g�|	'�Ԧ�T#�dݴ<�s&�D�ƺo�����IAH�r7�5�5�6�B�Ū݇��n�>V���bw�����L���Hy]���T#��V"V�!}V&(9��I�#�p���}@�]�Ҫ��F�/;v:�� SL����C�E�C�I��X}&F=�L�:Eژ��ӛ���+�w�kB���Ę2�Au�ر�E\;8F6*| <�:'v*�j���
5�l�4�ߢ���#"���8>/=1���F�����8���'q���V?z��a�K���6n�ܱ-Б-�5c�K�m����ma��1������6����պo��b�|/D���ӛ�dUiۤ�����*6�1�8���Y�x�+��U�y�LK�rw���{{Z@�3���k�bv���7ꑳ�����%cT�9�Y�Q8V�AZ��1����<�����z���.b1Z��K�f�A�ًRP����� �z:F����,#������D�Y@ -u[ -�G�G��f��0&	�s�Ĥ)�����N~��][���!�nH0a:H��0�~h��|���&�T-6�1p�%�r������N�+����T��ZN���%��69�"����qޣ3.fk�7���':�i�� �g��9r�y�}�d��|�ќ?�D�#yH%��$��g,uyq�H0�2���Tum�ox,������=.�66UՊ΂�������0S ;�vw�V�c�À�t�}nBź�)�~(���zm�~�ϧÇ�i>���n�X��?�=�DK��=����D�`����n�O���O�s�O��S�� ��qd�n�8娐�]aal6JR�C����8�8.��WLWj����qS<qt.iHȡ%{���� 5������j(�����)�#��R��_w5i@�l�W^'���L޽�,��se��;�Pdi����l�84J��ݟ�n�u���߀�Wd��J���&�����aƵ��IZ�,����lJ��M�8��h���*��ˁm��j�J�m������T�~�wƹzjL� ��v��0}�;?Hw--xDDQ�p���jºJR	�m�.���V��`ˁ1սE�ƌʅ����!��� P��Z�W�M|�}}uZ��ҶA?�����;�L�{J��ô`l��R��ᎪQZ��9�7�\YN��]��z�Kd�7��q�s���n���-A�����t���0!1FEN��V��bYb�����̥���f|�8�,%��?�߀	M_N'S�;��~�@�L���p1@���y1��1�k�u�E֗��7�2���ם���\7L�*�;4�nB{����u���0�� ����`j�"'��lmM���v7���:5����nn��A<2X���p���)2�4'��ؠ�bw�O�7��"���Nt|O�����y���cl	���W'ɀ�$UN�}�xg�{,�I����e{؛����e[#��5�T/o�i���~���mE �nM�0��RNY.l3q�ޟj`�ks6��U�R�D��y����ɚ������;��=Ʋ���� X�f�kc��&����s�6��)��Z��_�q洸�O��Y��tNZ�C�QvTm>1���L4��]�,�c!1W�d����G �8��4�}�h#Î��y�M��L�Tbև°\(%�O9O�f(?W�U	&�$0������y2���a�V�[���iLd�{���y"�a��>����l>��Qu�rB�k)fi�1r��]��m����_��1Z���d맿[�-�o�	��G��9���6o���u��9��u���Qi��6�:�%�p���X��X	��G��l�:)���56��iNm̅�aSpP��&Y�����W��:�me�iTO�O���Dc`�s&��4ZM]��^�M8��,����#���B�Ŕ�U�����h���+;R����b�	�S<����S,*߶�	�b2Cj|���"C�"@�衎!Q����~R���c�� Gl;�,#�ơ�-%X̛��� u�a���A�P≢�Wl�1m��Fk8�kꘖR�h�l�u?��Ꙫ��0���$�'o����sM�T�"�3/K�w-��&�l��Hc��N�<dGG��(���4�c�fz}�#�DƑ�b4{Ź�@|*�tsD��^0�����D�m���U<�ei���:�N7~jT��&�v�l��V�G@d�!v7���V��no�`���մ9h�#�Rj��:+���x��r�������L�u�����H�_��fd��c�w��:����9�W�"��F��v����x���!�X	,���G��s�Q��\����$�(,�������	��E#^[,����y�n�+���{�N�q���	]н0Ѧ���'@����5@�K���Ԍ�򣻝�y6��Ud'���L�4�_�I�6�T�H�GS��ޓ��dAj����Ɍy ���^Lw�Sk�E��u���(-���PG_\�c@5N�y��T�"!�^�R��{9P\27�� �%���Oa@��dRT�T��Yu�Qy|-5T����^/�ncuc����:�~ʙd�T9!y��o 	��M�J��P�G�p�I��י����kg��l;6Y�Y�hc�� 7jc6�@b��N��"��=�(���,3II�:!a�d�6L�Ʃ�6]1�*͗�S@!0�RI	�lJa�C��6#��x���ڶ�vWLmg�"/2(*�`�fo�λ.]s.�+1�NS�I6��	���2,I�1�h?h/�Fɸ���z�a53KW�
w��S ڪ��w6��Dj��Cg�$�ǹ�(N�ͯ↹�X��H ȏb��~�����v��u]J��?�*mb�*&{t��^�$p�VY�`��Z�D�����b������<1��%&��6h�+��v�?-x�*�$�� $��U�G6&�������ƍէbH���3�4?LJ,����nm��q#����z�<���
�����&B"'��D��F-7H��\e
���2[�,4����&��M�I���d�8R������h��_m�ڦ���^6,˄@�͗,�n'�D�*�=��k�����{�`�f�I����7Y�o3�x�v�!&s|G
S��<���B,�?��3d��gu�z�h#�_���:�NZ�׹w���JA@W�����>K�M�%��
LU�ak#[� .����� ��w&^d���=:n#~8FDD�SL�j�蠋�(͙b�e_>��5���I [6��p,��H�3l�d`r="s�Y*dN L�4��Q5�P� �؄��I�	��� ��-�6L:�L�w|'���7\�"N��p4L+���F���~�9'@��.ʄ�D1e�@�M�K��X4nr-T�`_�җza ���}��.�X\1uV���e��JX����[4	ިsҘt<>���Ÿ��Q�:�d
�\ �.TfpV�g�b�d4���"�o��!���Wm�x�0Pi�k�Gg��c�7�=\{z�ؘ��y�s�u���=�s/< �c����a�3�换�:HsUx	?%^H�V�39͢SL�}�*Tx��N��<����Jh��s����ў}$[�Q�E��A����V�v�C!:y�J�W(B!���Nm@a��%���4�Rf�n�*�Z)��i4��J��:9i���������q�ur4=;�A,+���B̈�&#���ﴝ[�ʄe��is��U�?�J�߰c�븬IՕQE?��MI�`*�I �P��1D��K/ubI�a�tyw��D��l�3��n�U���$g��];��Wz�>҃I��Z찡,)����{ 'L��Efx��� .��2/MX�z�!�uW�ut8Z�{Ǟ����]w���;��{�ңO�(T�~;�,�n�u�����Jc��Ļ9���F�cˈŗ2�N�5OS&��6�2��#�i�c�� <�@���vO&��?��k�d���Yp��}əyUO�j�I��[͊��ȅy��h�P���Z��<g͑���y�g�bF���h�����o����J�D/��H)�C��h���Ѱ�.l�wsrVd�J�&�nl��=ת��Z�s�x�Ɠ��̩����9/SN��Uk"th{�u`*�L�2���O�y���[a͋��U�pL̐����Dm�\1��_��w�t���������Z_҆b�r��A�=+��Z�� ^1t�h�`@͹�.�@ c�f�TS�r�0�tSD��9>�E>���M�|�3��=P_m�5Z�|I��7`̀0�O�yL1)�T�0��"���?�gΆaҔ���=��H=y��$i��E����4�>9��(��=lz�!��*wZ��o�!��p=3٢�馆9:[�x�*兺�i�ôL�1��U5%�yO宭~a�gp��r1�ln�Vؽa��k���4*5�M6�Ϯ#^��mA-nsU������_��X ������<�)Ô]8�T#@�TN�p1�-�-^S}	=�y#:��(�I��n��U$f�Ţ3�OF4U�m����ǐ�-�*�2w4n
[���A���u��l�{v$x����Mc������8�Ԧ(%R�b�k�-ΐ�F���A>��Κ���[�>'��aqi0��5�}�vHEgf4G��(��C�x�|T�b�v����e���$�b��4� �8h֊?���PR�PÆa�M�UeF�b�0:α5�t��b���Ƕ���~���'x㼃��E�쓣�ǐ4�i����dw�_��88�q��ȯMHf�O��O��O{K$���o}�mx&�caC>�M��lBm��ZJÜ=t�9��A��p}H)�4 �L���Z��rvR�+��xQϣ&(�C���c4��{�v���fZ����V�@?,�P6�ҍq���߇+[���C�l�~.�B��}u��3���������>�q��w ٰ��qb�E�K��\�8T�W�P�{bќ�؊�@o+O�l�1ck�sN��b�v14��u v�k�|���Mm �JP����t�N�mJ�FR2�χ�r��gK�� ����p�M�����][O%�b>�u_�y��.��i�y��z�F_4)�N*&����8}�C�|h��ƽ�&4X%��)�1��Nt�� b4�|��^�����p�~t\WK#=?٤�7&X0X��7qM�u�>��P��z���1Os��ԛ#tA�ⰝB͑(\<,��y�*Oi�Ǎ�k�j`�H!l��^{�Ԇ, M2��t�M�]�~x�9������l;}�:JٹAhW�υػ�4�:����g>5��{G�G�Ɣ���{�d�pZ�i���M@�Q{Y�\�,|�(h�-��>s�b`@oB��!7�`�@-�i��ձ�w��;M�[�2�����0}�4�Ʈ��Թ��&�'`�)�h�ąцmdJ�7�i�;�e�.�5=�6�!j��LE��:�1BE�]�o/�dX<�;�V�X��~���u-mm��[�&p�K폩�*D�cE�m��+�q����?��7��j���E�:��8�4�ά��-�e�6F�`~�F��ɨ㭳&�OxM�Í�!��J�]T�L}e'������\rI��)4�̚��[Qsh�6�����g�"Lt�A�mW�;���zo��]s��*�$����7�ɳQv&Z4ׇ)��DS���ֱ�U)�s�q�O%���\7?u}�R�� <��~2�Z���:�m�V�7~��n�X0�{eI��#�M�D %)�lXn
�D-X&]]
����w�ˁV=Q#x0������XY�9��`?���A�Bw2ؠz\|�%�=g�Vb`���8�(�R�6�Z�,�(|�0?�[��f���+uw��g_l����R���{�t]=����h���͹�ۻq��c9u�=?-����Ѐ����f�O�A�T6��}C��{��k!=ɀڱ֣*RZڶ-]x��q�\<5GD�AJ���j�ʆ�EK�L,p��DV�A,3o��*'�5�x���4�bW}Ւ����2���lLE���)�)�9�Z[јp:M�a^����0�8x8��ƺn�ޝvM��R�J��봲dp��!���j��!�y�!��`�~O|�h9USv�����bP�<7��s[�;}/o߾��J��P��CM �φ=�e���w<CRp���ɚ� �u�z�f�Bz<D: ���������V�4�V��4�;�U�
J�z.:c7v��b+u����\�zt���+��Jm@= �/�ls���NX�ֆgp\�6R�̓��IT,#���>,���<�y@[�^�p��|�/-m706)l��ǾKҒTɲv@��L�(;�_�C<�t[&�!5aOEV7�\%�fٔ�d3Un��̮I��,L��t�������Ҏ��Vnj ���������Â�ۢ<�p�2F�X�=����x�׆�g_�3�k�N[-�_Ӊ/�_a��h<��zի������b��y	��M����Ǝ���Ƹ���Pg-q<�1�VD��Ą�cFN�R���ņqİ�c#�����H@�{�1���Z��G>��gs}#�B�S���0��t�B����4�)��ͼ�YX`���d��VǦA��)�dߙ�����wsY�����&��h�Mh�^g*���2�u��D��J��##b4J�d���W�WݎKQ|��F�_��z/��)Z6m������1fz�&�+�w;R���=�*�T���(�6����i �Q�����������t"7�»g�]�*[1�JЈ�|���&��;y��E�Z4f����/��/��U�w��Ƅ�������Ռ��,:�x��Ԅ����,7�gΑt���"�D�v�q�^�d�n"�5^��].�=u�Q�%z�SVY�,M&j^�E� ]4@g�k��t���Rw����NZ$��>O�:�l#;����a��`�k%{��D����dV�K�7�ܤeD#�Q�����%&u;Y!F>�ϭ��ܡ�c$�W��@�k�@�=8f��d���	��O#�@��Z��f�H��/��<�ǔ�̟}so�L��\J��d�x�4�Uڜ�:�����»/ w����S�{� �N�O�7\�%��漺c	ӹ��8��8����@�<�W����^���?�A�|���p
 g)�J �u��i�J�H��	��c��M�O�9"�BMg1��`��6��K</�=n�Ȣ�jL,�E����t^}��n7��G?�̤��o�V��?�c�H&Z^q��F�͖6=���m(*�Ԩx9�l����u9�B�<C�3����^쎿�|�QAP|��i����g����,?t���qӪi�X�r��QZ�.�=,�Н��۲�86�3�̞�&4������o9K�Öp�=*\P�|�|%�E:̋z���Q���'A�.�.��-��R��[�/�4�yf�h���%tt_ڴ�L�:�K�����I�'w8I�X�g7�����L�Ns�\�C�x�.,j~ǃړ��o�Zݸ���x��,}��ż +��a�~����{i�<G�V�g�o���-F��GX���7�A�LII�-;'t�Gi�9�	kZq�ZZ,9 ��Yeɟ���1�ͅS�6Bm\&P^c��̚�����o~�g�D'���
��^���ڧ,A�h�K]z��=�n�s�$%�Λ(;U&I��p��w�kE�Ջ��zS��'^���v!��n���t�Ъ�g��Toq�$�&�y��=���-��>��1Eԓ���H���~�k���yc��s��`S���v��
��9ڀ�F�^�"�g9/�}���ϫ�ql
ӈ�&��)}?ޫ�RM;?�Fvg�����L$��g�M�lM�����{W���4(�Q�m���A�Q&lQi���%��}ዼ�e� �o�,�ʠ"����4qq��1&Ј!�Mws����C��uߟ]ߺήڻ�34���tU�}���~��o�L�͂�e���%�}w�Y�l���#�_�ş�m=?� ����;�JzH:nS^�G��f��m���꺧e��X@��>T�	��I}j=��'�i�K� F�*�[K�1.�H�"`�#�=�;-��Ս�S� �7/��J9�tL�]�=���:���j��h���§�?��W}�W����� �l���=Z�a-�*b�����P��А�I9o�sp�3$C���%v�9
6j���YHK�cx�+W�){�=��ǚw���}�io�:d��VN1a�ӈ?����5f1-J� ��u}�����8�1�ڎ\�1tP�k���ph�f���h߻`r< ����1����ZF�����@�7�ɧ���y��9�G�gl-{+4q��x�w���K�?�5l#)	��d���7�Q_����m~�����?�áF� �����-�j�Z�	�3��w�l
�E1�Fx~�NjEc*�S-�������,�������(�n�A�,�n�<�ƪC������,�^���?��r�1�1�a���@��k0�<c<�}A0�LdDk"c��D�0��5�yM�,Lt�-��|�:9��ps���
/ԍ{���%�s\ �L���߫s1�k�ZM��v�=���:4�|��=~m�	>�ȣ}Vނ��*am�o�$(����� ]��DR@ee�עд��L���M��s->��S��a�Vh߸�bΥ�+�@�i�V�㈾w��L&�X��|&�'�-:����8z�� k�ױ��(���h�=Jm�[�='������c��1]ڥ�}%������������gǏ�e���0�X�H��������{��җ�z׻�W��U��^����BQ��:��g:o���q�d$�ϩf�!��x.��|��h<����Ɂ�s� �O&7�a�j���y��"i�9}�>�:4a&:x��v�=��=%���:xC��?���q�1ji��'e<�$��j���>��p��Ӳ�r;l�9��F�h?�X�z��Ds�-?WP���1Y��QےSЄ�x�䕽�g���|ڧ/O�>;oww�L�@Ts��#uw<�Q8�_�K�z�C���!L���.��km���\�7kx$Ր���i���uԴV�D25�!�$�M(��Arۚ�j��&9�右ԧ��&��Y=����ܝ%�G�8Q4Kj��К�h�Mb	UcK���I��Ej�q���ӂ�j�7^?S���}
D� �l�%�@t�l��؏�N;���4��x��;�A��a�CA
l:�Zt 7@ȿ����1�wc���xy��έ�,+?QeNy:W�T��A����tB~��4#t��9�����P L:~��++�k�d��%l��󶯐F=��bҁl7q;�q�N��ϊ�eT��+�Ep��{�찱h{��h(�Px{�U��bqXwb~Ѓ<�=�Bq��;��Z��p�l�V��ս�����xf�+����o�����u2�E�䲬e򢂗א����w�m�L��woHmE���JE$�;񼎜5���j��<���g֒�s���¡W^��J��h�v�ԕ�;�I*�}��M�����1�<w69���4ۏ����;/}�{1�q�!�`�h/�%�W��v��3t��*<�5nҿ`�t�%T	 0A,���J��i��dMx��Tc;+� �^F�X|�+^Z �����b��H��9��z�iDB=hh�uZ�	!��M�T8a7_t���/���MozS�����z����LQ��jٞ�w^=婟��M�>O~��.���uZ�b�M�	�ޏ�&͕�I�����.�&<޽��~0j�ߠ@_�}���{�Gy��j�m8]�:���e �յ� �~}/�����ﷇ%���b*�e*m��LV�{�}�V�Ϭe�����;�ɽ�N����'}��<n������9�M�-"���֠u/4�3�o����MGM}LD�g�g���~پe�|���򓰧r���w�^	��G.<�>f��$�>j�_��=Kz/�˒����0w�F }��8yv��P�x���ȏ�HyBW��ۿ�` �,kS���Ll8�+�`]�h�j����x�Mr��K1}����i�l��F�0Ԉ��-@�p�7m>��Z��08՜h :�����9�A�\(4��_X.╯|e�v��_����Mf��|�ה8a�w�աL�t�!�Xj�P���o/IT�"�c���"���m����H����E��P���nF��{:��4�+�t��Wڍ{Q�`^���)4���1ͥ���̛e�qn��/[��2Z�N�^��j_d/~��/9m�� HH�0�8��YZ��I�i�b�2��h!3�.�k���~˷|KI�b�������_����q���Z�8H0#����#iK5^1�s��(�;ڊks'�:���S1h/<:�4��0�c6�/� �0�y_�З �f��	W���X���r�(/��hDk ���[�Z8 �6�5X�h ��6���P4�-����/�i�&&G8/N%TƗ6���(lo�y��h;�Q��+���ލY��P�	J�ٞ;�5�5����.٨�[����KS��C�:�/��m~����e;�Ns�C�oM#��VǶ��9�~��eJM�b;-@���D�Mjg���?�Lk��U����#:ɚ�ʦt�?������</Z1|1QS�IF�Xl�yL�.�n�������n�c���h���~���Hџ�n'eXSDK��~o�-��xz�9�yn����U@5�Qn�tP�����AepM�BY�$�O�tb%b�"&��m(�#@�Fռ���a֧E\�(�X�Nh�=G�$��L�}�Jj�Bo�8�+�X�o/i�MS2�F@_�z_�1&K��q��@g5,%��k��6j���tr&��[ṿ��9���~n�:�l���f���f��c���|�*R�s���T�N��:�Rt�3��"qȓ���F�3?�3P���"w�A��:d���2��5f�N��҅k��v"<ҡ�mw��s�E���������~��>�O%��s��9�QXa0G [�4n�B^����ĺA��q6�f�GkF[��a��m���Ȟ�zm���J�-��1��b����%;���(�4����h�.�6�������<���L����G�5ړ&�0Q۾OF��IC�)��t�3�U[�di� �����'�(J���SN��c\>�
Se�c3U=��{�iE��v)/���X�k��et�d�&< #��%��ǝI������'A��zqqʸ��X|뫨����v����%�΃a
�����8P��z��Zx`V!~Ҙ��h��2��f<� �f�3L��c���Vɧ���������a:��߸D?L�^�-�/��{p�H�f<�U���z�Rf���Jv�25rѧ1�b'[)������Ak�{�5C�E/�C�r���]0�H)�v Ϊ���d6��A�+�*C���=L����0�Z6Q��M��K��,������OxN�b@�H�YZ��BQ���8���F�P�_��Хh�p��x$Z�֋�#JC���fm���a��br��,$�y(��)��B�~���8��|�s�j���%����3�+�n���9�`8�㏼[֝��u��M�މ
)��P����Ė�:g}�>�3���[�Þq�E30l pI�q�ŰS�
����WO϶��%p�=]X�e���	_�����r+���Y#�qյ������I**���T��SW[q�G�s�	̂ߑ���6�Ęm~�������6܏W��CJ��35�<��qԁY`ֹ�9m`Gٔo���C�?�UN����S�=�Gn�r�͵�5�>�f���2n@$�U�m�����0����
���Y�*��*H��Kj���gL�I���Jl!�����"��+�q��Җl4����Í�q6lٛ��sQ6U,!-�i�ϕKI�a)�c�5��4SգNЧ�r���;��>{Ϻ�p��!eF=���xnk�x�*ǷU��T��y�kA����P\�7>��ris�NI�	E�@;�O���	 ��9��g֥���!:��5�����3�#�d�C�ס�}`�:�Ǉ�qR+u�T���d�)rKj�5a.@g���l��$鷋�,'ʃ�ڎx����)1F?��	���5{V"ߢY2��t�O;-{�!fK(��]a�rl��#�mn�܉�o�yE����cW�����)��sM',�4ڥr��γ�x�JTt�o�(��Ӷ=ǳH�Ů�N^��]^:��c�T��������q��,0�K�?��w̝Sr�����>I��G�N<��?h�y+��ޠ�V�w+�![�崒���~�ߗ-���4��΢m6�|: �z�W�M+<����V����!u�S�~����I
�I�$��5g�4��ٖ���rF	̫�n���~�����RGc(�FU��~��wV�
M�,@|r����b#�$ d~.�m�(���滕�|��y�vS��*�=��׶�x�ss���5�+	���^u����oAz+[yb�y��e�����d�9�xf^8#�ڱ�f�me+[�����8+�x֬R7Q/R��i7�};�3k�.�q���)�-'���<qe�OhU�^�y���*���	�N���n)H1ۛ���>{��|�Q!q�f�el^Vg2hN��5Ӕ���6_�Xd�#��B��4P���m�t[9��s|���*ӯ�`�
�O9)�,���DZ�s���\r��N�:���C$�`��kȝFΛ�h�� �i��I0�9��w�sS�3� 3��td��c�M�����='\J<��O��Mg����+[���zG1���������9��[X�
jf�X@�x�6�ŧ�\�L��CLY��j9S\�	�)'i%�����}c�yN�e�b{�k�Tw��϶V�v�=�ռ2=xUM�z�;	\3�vG#Y��y���!�o��3=9ے���Z�s/::��r����ֿ1}��`�G��Ӿ�uuz�v�;Z�԰�O�[Y�F��Ew�����+��Ȁ��C�bn��dCԓ��6<�n���f�]F_�
���� |�y�8�:���R�:�cV�����LA��%�]�o�9ۮ��vzזF��*P>�O�`O3vΫIg�Zֵ3����cb�J ���Z�f蚒L:��ӁUVU�������pV���R�٨�����bSv�����G�8_W��Q`��Ǽ8`�N�!_���`�bd�d�[�˕�MZ��t�ֳ��|�C*�������x��ǣ�2)kJ�,�L9	���]{�8�D�ʸr��IB�����.I�X��8z'���ˤiR����u�[��B��Y��ZH���w05]��������(u#����N�v
��W�."�[*3ۚ����|:m�����H���~g�8ǻe��g?��e�^��GTw&
�%.)�p��=��x�41�G�����5A�/��//�Q9�FB԰���J/�&���i��d�{M7�,̀��Ȫ���4A}N~2���� �-s�%�U�A`�
��֝+�iL�֌�ɂBtn�$����Os�ӊ��|/bXn>�q�VV������g�
l�6�#���T��d&xC�]�Q��1�����e8�vvڡ:P�}4�\L�|v���^���y����BV%�C�MHV6��8jx��g�8��]3���W}U���5��k_�ڢU��~o���		`#TB�o�x�UZh=iO#5�X�l^7�s���6Wq��-w��=��K��w�d?���bCaj�J��~�p.B�c�t�*Mv��c>�Rp�0U�jk�*��Ɗ��������+|��e��?��?-@��(s�-Q��������F��=�tI�mt� ��؎x6���lY������K��-���4��<�J���'�̆}��^_Zg���AL�p}@͘	)���v�s<��NnX����ҳR�9�4�yMM��4�$�z^:��kgIĴ�r���E0�m2��ww�I�Y�d����}�Y7�Wi�g�\��������h��'4�t�%��ri�_6��P��$:��������= �`}s}�oJ��:}Ԧi.A��Jw�	�N�CǰR����̧����R�݊���N�Gx94TL^��/yg7
u ������-��_�x�7U�9���lYM#
�4$�cʥu���x��G�e�H~�����owQ�3��e��ŹG���zCG�Pw����7�U���w����y�i�o�9_;p�x�\���_�=��X��F�<Q����;w���j�75Ԛ�Y5�7q��ǿ�����:Kd�Eܟ��`Q� N4Y6����_��%�HG����Х/y�K��P����(vL>�x�q�A��<�X�+��+E�ĺ�6�:B)��s�^��3>�h�t�������_~xٱ5#��/�Ơ4 Z1+��ԅQ���c?�cE�������5�{<q,�����tXzVW˨�ض~���ge�N6�/v�M7GlY��Lg��рp���-F]�-��>�V�)\^S�zQ6���iL���x���	��l�Xn�Yvʘ \��&`s�L�Fv�6�^�ٕ��b���^�κw=�w��)�=Yx�S��;C��E
�!���G������@�����.)8:X\��?s˘�l�c��������n�)~�J.()�$�%�[K_���
YJV%��5��?�3N_��]m�F��>�s��������׽��2�%�k�7ύs�x�[�R��s"`;%���/,�g�b ���MHݐ�cxfϷP<�>�_��]��3�\��~Y��\h/l��áŲ
 �L4M*�&C9�2��5�8��b�¯Q�cJ�-G�dr}���+t�7}�7�p�n� ��|���>�w��Ґ��W���/;-�^5;��y7��zf���x/'��k�:��4�vV��Ѽ�9[܏5�3-G�_]�X���w�����~��q�i�������4%���]:&�Bq��N��?[.<�fm�N���:ۦ��6�� yw^0i�]m������,���e���a�q������������rZ: )!��DY�?���B�o��ļ���6E����j�*HI
RF%����J:�yf3}���v'�|n2̎���:Z���Ԏ�Fay=#r�C��ъѦ�+�jX���.8N��\�F���<��4�м���备?��惥G�4�<
/�>N��4.Z1�n��G�����ſ�e C�9\�E�x��ye�i�@��݃י���ʻ;�d0�H�{������®C
p��8��i�N#�ǃ���Ԇ���>���]���+�9$â�@��]>��� �N[���f��כ��N���V�!C����u�$w8N� Iڒ����zf,��Ay5n5����C���h�Z��|9�w�n��N���]��M~ү�- @�~B����]m��=5������:��J8�981g9�t�����__@���/��|M�������=yN�%�{��9p���X&�:F3��4�
$44(N:�o�UЇ�@�pV�*؁�����}ۣ�f��~gRUx���ܣ*�s�Hh��X=��̎1\�kp]V#���X�8����1���t��_G��L�N�m��k
p�A�l� �u���ɴy���Y����On��>�\��)��J:�n4���f�j7h�,�\2ل�/FJۃ��M���#�8��a��Y�ni�䈻����W��z������>�i��d�e���Q;�l�KS���a�8q���1��d2��kq}���o~s1ɐ�]l�@r�����jS9/X��"�����T�k5U�Ѽ��C&@e�WF� �=�P���8)#��r���� ����/��������.�>	@73��*����:�ZY����H�r/>�	^l����k�q~�tD{p�i��Og�x0CC�/������;�Q��2H���n�t�����1��A�P��4���e8��t�<�q�7���{�o���sԻ��2{��g~O����o?e�\ߟ�ĕѸ{����f|�����|�k˅����\�
�:�����y8f6�μt굝	����{�m���zj��]��|b7Jz���μ���Kʹ�׉Tm�֜焳�4����O�����51�c�#�a0�%���ó�w�$}PG�lz�����ڣs�߇
�o�D5��\t�Ч(C��I"R�ab���y<������*��+^�l�5쳨ȩ4�ǻ�#r^h�!�ͻo���B�uhC���]��`ؓ������9�;�Q�K���R3���0$)�U5	����1܄I���te��il&4�<&/��{L��FE�̣%��	Z`�v���9�yN�_���=�����z3z�Ϛ��?Ҍ��E���pʝ�v����f�x������
���9��X��ۚ���m�#�q���'\9����֠8=:�|��<���7~����4���;��4�?��?o��)f%m�IY:w�(�3j:Vs#VM����F�߹�2�є�������KG��[%O$�w���]k-��P0���
���j&5���� �;ᤖ�xp14�
�bFF�E��TԸ4�O��O���~&�@�@�p���Nk�q(�߶�J���f������E;���bAx4���X�i�H]t���<��Qr�#�K�A�5	��������w���~�����?����K�S*��iY'�����9ٽ����a�했("��rOs���6�Gn�kݽ;P�>�5�����DUtϰ�<@�eA <��jċA��y	q[ x 7j������aG��l��~�fr��4�w�^�R�_���i͍eȽ�������Ȣf�+>����t�jN�vP�Ŕ�İEǄ|�� ��2՟���Q󹧑�4��,�e�8F�4�Ȑ6R���<4f�B���!�.s�����G ����/�Ғc���1>0V����x�:qG�v<�� 	��ul6b� )�����ީCv�"�l�ߘ  ~ʻ�1���^}7�19'AY`�U�@t�\��d�!�|��w,S��\jr3��t���u2��Y�o�3��/�� 1�~���^������ ݶOp��xgtown�M8*�o7�G�zFɹ�l �f;*�C���#����>�eQ����B��17�g%�n�so�'�EHl7��t��$����7�a餱�\��\fB��aB�w<�a3�ԈV�9�<��"��1�E��v7X:!���Z�GbÛ���%ݘ�ٱ.06���s�S�����^FE1f�d�b)�S
��/@C���q�w͒��J�»�1,0\K�� ~1�LfW�y��� 'k����d�3o��t��:�lR��S�0'���,1�K%�a#����?��������z����^wa�&�>�w��J�/��Bw��x�1��]�7ˊT��g���g�����w�%��j^��� ��r/�'
1�=�)�c\�3F��YF%ԭ�u�6m�{���[!�#�5^:2U9��s%�ΏԞ3�že ¶sj`ϛ2�uKԚ`>_~��+�4<FM/#C|��}k��e��mb"�����$ţ�{ؖiu�����?#e��/���:���A4M�gU�}��h����3�5h������0�B!��+�����@�ö3x�;�b��h��ۖb�c���}�� x����m��ѓ.<Dmr�8�;X��$n�JD�X�G͠�l��>��lP^NS�I׃�Q��`p_��t�f��zp��C4K ��d-�bH�P�1�GC�D[�[��-l.\-q��$`bu�
�nw1-�=��Ym��g[��ܩ@k�Q�f��iw���s��<���!�u1x��>����Ӄ��6?�aT��}n�V*����i�_��q�#�E���J�vҪ��g�#Z�z��D�tg�*��E��`	��o����A{BG��K��E*p����g|�gM8�\�
k���f��Nx�N�����r]�cn<A�;L����ދ�[̎�����w}������9 �%-�����< �/%���h��?���+_�ʢ��Rq-@��~��=Scs�_k�7=1j+�K�r���d��~���Ƕ2�Ƌ���
��
`��j��<˵����h�]sZ4�/S��� �{���(��gy�����֦2ʡ�`yέ�'����9c�gE) ԰���ӌ�Ur+�?�Ll���m>Ǚ��l2l*��N�U��E��!dFڀ�mԎ���}3]�������Ԍ2�j�M*�:8j��j��1��.)��������F�x&�{��dg������ާ�|��|�ou��e
1�B�X�,i�j~��p�,��j���� M� �C?�C%<��D
3�S���?��'&+�I.����h5��w��.�5��:Zby��?�Utџ�����= ����pˍo���FK���g�9�3�-����V���)�j�L��0I�0.+��>�����2Y�{�[f*I� �IOhp�s3��J��#�����7��lG�-?����׼�5K��Tz���$�E>���b�
m��m��K��xi�Y���+~r="��{ǳ.(tp�4���`��J�7�s�< �����JQ�?���^^Ƽr�L�/����g�'�Ά�g��w<�@�Ώ���7�����*����'xȐ�*���w��;���4���}t�'W,O�TKr܈$��YIY��~�k�,i�vI9\�p�����V�yQ�0�?�5�^ĤP$8�F�q�d��i*譺f�}�l�xUƁ�pnJXg�7&ΝP�Ƕu�:�y'	tL���	��.�i��iZ�e�#ڌE���T�Q;�ְ�KL��{<�[) ��Ǳҡ*����^F���3��+��F�ʚe��D�v�],/�;�|6o{p$	bV�B�������i�����?�3������0�LWE g'?\ +�8mM�7�́�F��1:�t��y���=�I��a�mh�ĴP��輈�y�c���%h���+�2_�K�`1���G��iz�F^*��c_��p��w=o��%�2g{�U��YD��@ƕcV�ؕ�BVQ(�~�v�"�P;M�0��a��t��r����n�\f;�FX9?�#?��Ji)��:pI2L�V	�i��*��H��b�p�n@��P���Ң�br��Rk5ᲂ�g���U��'�������_�P���P�`i9�\�T^���2��5Ip'�k1>��P{p��1=���P���0��h���6�`�4�u��VJ`t�`;4�v��zƢ��h{��}�"F٠�>zTz3���db��n�i�7�V�!�b�!�����k�.�L�̶\�ӆN���r�]@�	�x31�	Ř�B2�`���w9���y����`&�P@m �$�[�p�EN���#���a�o��9���7\.r\��W�W˸�^
T�b����厵��� l��.#��;�]�c��e��y�}�����>�++�����e/{�T*��@+f�#�5	-�jD4*�5M��#�w������YrţXƲ!���@j�\S����'��m��?��&R�?��m9���<�v(WIŴ�a�ʦ]�UTø���7:R؇�rM��x`GM���M�0T�,��5�=���Ti��J{���&0ƨ+�1� �L@��z�s�*mRJD�L��ա���=���y�UϙV���z��h�EΒ���������^�e,o0j���Z�]�\kP��0���;w}�8��Y~�t��MтKxǨo�v�.+&B!Z.��I%�C��$�����,�+\H4�����E����y�M��AZ���k��f�[��҇�;)tA���i-��I���P����n 1�;]��d�,
1Q�<�9�z�C��@It`M4J���I�i�w�.f;��Ш5a�n�!:�se\i�}e�{��P����Y�6��&xL:�,���P�K>O�}���j�h�W��ssFDʂ�c��]ES\6�՚�����3ӄ��p���3���W��ʈ��s2c�3Q��Q{GjJ���Y��*|��M����琚�����UERyO�,������W�m@�O4_�MF�a�؋�D�Mmap�Z@֬~:I�^s���r׃�����Lh<9 ���@,�cxʺ�آq.�!6���>a���b�y�ա�X��N�^�>Ԫ�k��$�/�|�ŐI7/��6r�Ӿ�p�G[�|T�cvx�2�}�G�N�p��ֆ}������ߝ&m����;A;�]���7�H��5��^�]Ԑ�� 컬Ɩ ��S��[)����T) `�A)(O���ݖ9��Ox��ؾm��Eu��;��5�ub��2���;F��
E��ǭd��4G�z4�A�6v���vz�����]c��!"�-������_������DD�������DN��vI��(���J9���c�t�[-z��i��@� �7�םE�b���,i(5d;_��E�>L��:�Nt}
P�������n�?�9}bF��`::-ƣ��8�BS�`��{��y��OV����5̪y{-�L��_�М��:7�`x��]����&�f�qK6��k9p\�LS���˘�����s�H����0�����8w�ü�>�m�'_,�Ej�#�k��r�X����/[zxe4d۝Oh_i�:6�󜩮NNk	g(�f���]���4|Q-"'�I��z���8�?]�y��U�g���}e���6��� �S>��T�ѡej4
c�N	������ͱ�bg��eb���ye=�G��e��KIj�Y��Q�����V���gu(c.5r�F|9�etD�\��2�@O�i3�ޖ���%O��h��q��C��@Q4͐�Ԇ��o4oz�p^��#��Ϛ���y�� ���i�4��K��K�c5wK��S�`�������\��2�����bD�h��|&�F�  ����ʙv�K�#�A�I5O���%��s;~�0�q
�X3ƒ�ZL����bG��[�8VoV�<��c�;q(�����G�;��lMO{�\Zne�|ѓ<מ��6"W��I�ϲ�O��
7.�b���b��ˣ�~�i��Ѱ��臅9n�,5�a�m�.� \��aw�r���e��K9��n�䖘�8w�-)��I�֤SՍi[+ֹ����\��px��"��H� �n%�'��Lx�O+[ >*�Y��{���;� �Q�[��i����� d?�ղAT�tzѧZ�n��δ[!��!7"M��,؃�1���5�1��\k$�&b>hz�=n]�M6P6��D�"�^�,<}�dE�-o�Š�6�C���D%Tl�GD�FC��v	�}a���ۅm3�I'̇�����/'��B����$B�\��E�d}zɉd�~q�p���=�p�kE^��o��>���br͛>��p���b;�|2� 6����@�����������PD��!�v�����-�(��89�R���;u �R�����ùA��C��b'�\���4�hy'{�2jkz?3�z�j�E�[T�#��Eq�M�}�F�ѣ��0���Y�}�B�y�_Fß��S�-���:= ��5`�~���.�ğ]���xt�˄:ᤗ�#��0~�>����E�r�3���$9ae�o.�KI����n`�������Ҍ���Ck9�"�5zo�Ծ �D�Q	�BU���tgֵqLn��l���b�"�f�+�#��!�����q���06�Ś$r�ir���p���^ic�ϫ�,��y���5�d�<i�����}P
�+�޴_P�r����;ݻ�'���-�佾p�Z��� 0���$�� ��|?n�3 ��T�m�v�9�>�P}gҗ�$�����C�4�A�b�E� &���N��?G����wfJ�����H���=�f�<~����3�K��>w���,��E� ��O���L:�c����\�f�p�s�#<�� ba��n7�`cD����y�~�ﵵ[w9i��]>���Z�����T�<��r|��i!��>��n�	��^�e�|���yNrKZ�A���dY��6\�Or��4f�
�6bC��i/��ݝQ��b��w�"���?���w�u����'�3k^��Oo����ь�ԁ���p�0�@������=�KʳsQ6l�qGjMFG̗��)Q�W������/��Z�?|w��������,?������I��䈗V:F3�z2�u�s§s�<��wy��Z�~!��	��K��i{��/�}�jR�s7'�׺�%�!�Y�s�c	8�6|�½���IVpN���g_�&w�?�2+��"��$%j-T�uP)i8-��VM%N�M
"���m���ȉ <ߝ��	�1�o�C�Iz_Xo��v��m�Iǭ��Q�� ��: �
#y�cް��n4��N�8�s�\{��������']m���4�Ϛ��^�	�V�\����i���v��� O�uϸ�(�1!o	��.�Z�?$34��QҔ��4�����f1n�=6o����������h~Os��f�kÇo,9��l��� �@�X��Vk	�Y$E�:'�13��u�F���@.ԙݥFc���,j�	�j�����#�}e;Y�H:0����ZD�]�<�@&���t��/J�┅Z�BI�vͬ��\H|9Fe�s�1}&u�d�Ny��o���8!`6#'w4�!�)�|n��q������C0o4و	���`^���5���;�+��i�;�=�u <jw�G��7����o����G3��x�B�̺�8�+�;�3��<�#��֯Q�yo�1�='<ҟKi��W���qs}�j���,?�9���^�����Y?!M��:����	~5P����?3lP�H�tq�>Qs��djvu��<��J�El�s'H:�k�C���j�ׅlՂ��B���Ͽl˚]v�Q�~�����ĢTH�����\��K��9?Wj�w�B��4rr)˝���˻��VM�H��M �)���~q��d2e������}�}����
�ģ^����op��Bmt`�N̄�=>lf�Ǔ��mv�����G�R+�x1���f���
��;K�[,�s�{�f�=;��w�i����'�&��u��i�Bi��Y������8ps��䲉�����f� ��[J��Y���L�o|�hC��vI߇��{�+MZ�	5/�B�8 "��\�l�Զ��_��"Y�~��h��
㣎�Jg3�vG��K��M��']QYb��E�1�]�m�сK�7����M�aP���o����(�8�(��!	��,6y�^�]��i�;AH�k#S����D5L�;E��ܝ�N�j~v�Z�쀁Jڤ��N��G�C��I�7��l�[hD���yoëa^�O�JUƄ���3�#�ݻ�v�ּ[�g���M:�e��B�Lk0犝INZE
iS�\���F�Ms�|�n��H�I�$i 5�z�y-a?�HB��%��\���+;�����.�%�8�|������9fy��M�q�9�.�i���RY�]��x_����N�����H*��?Z�Z�\�S��R舝����qK��x�����g>�����MG� ��>��>�������	���Ex�z��M��'�w�]5����گ����4�ɚp�{s;'S��` D�:��o�S���v]с!pg�u�2��R�� x��h�B;�Hs���=�Kl_�lT���;*�w���I�N�E����vJ!z��I� s2���}վV��&�hN��$Qp��U�e���,���_u����[m�;��&X�;��L3������,�z7��zK:�8���g�{g�*��R�|�צ���5��`{�Qv����tW�a��S`?���
ճ�/���M�E{r 2�a}��=�䗣�R��偭t�dc0�͢!�E5/F�d@���|��k�v�-��}ٗ5�����R��S>�S������y�4���I�pߑ�i��'�)`6kv�t����$:���������6����N3ݙ���ʼb�K�q�媜7m{_簟sS�B�m�
�/F%�uP�.��,�:��R�S���2���a����i5��&D��I-+��UϷ�=]Xұ�.���;%A�62�$�$���~�Gf昚r}Q�I��#>na8�����pQ�8����He����X��۫�i����2�aB�)�d�L�y>nK����fo:��N;\4����m^���u ���D@��Q��t�uP�	UbB+6p�m�8��������������rr��. �M�m���B�,��Yq��Wq���i�;m�A7�4�����.���%��D�ᜦ�{�-���=M�h�(�[�7���^���34��B�L���g���M�U��i��U��8`O0������o}�Ȫw�%��:�v��V����,���*Kc���m׋��'}?��Ԁ��s�����)��җ����H��,T�wql��
�DBsF�d�$wJ�e��%DGt��|>k�by���^3� Z(+����̔!�A�3�*������AU��N��1Qu��hK/1�x��P���_~SQo���Tۏ��ਜ�j����̫�O�����Ng�����o~�E{���[��:��;P������������%�4U�<`	8���;8������B�4I*ƶ'u�Be����hĀ1��IB�B	g]xNք��j��3�ǣ^�EM�Q��}������=
Ʈ0�4B��3xd�EB�&�AS)�J�~��_] �M���Ƨ1�\f�1u���[��ǻH=AIRnոv�/���7��^���BD��C��98� p��Z�d�ִ�����hJ?�B*��	㬫�
�ˠ#��a��rŸq�F���o��  �8IDAT<�Tf"ځm���0��[���#�#<�+�u�t�����7���s@@������r�g}�g-CI|�4�.#Tf+[�ʭ*��|�(k�����1��~�`8b(���~"�=h8l`�N��p��ɗ�;:s,������I�LZ���7t2j�%=�{�:x �z�]@j;s��Y��Pb��N6VW>��>8����#/~�~��m8�ʩI������l�NK ��(���r��}�k�e���5�w�,�T�����"�YsM}N��3�;P�4_��k ��U�$�����9��\x�p;u�(���7��~�}�'�:�������Yіm(x^�u�4@�W Z�i^�"����%������s�G�u��	��2ƶ������܇�D��bf�z6 _АZ��V
x�N˄��`����%�ŀ�5˥22�c�j ���,
���K��&��ɧ���-/��ݴ�_�E��G�kK\kF+���Z'"y�	�ѐ��Фx��^V��[���Y�X�X����7��7�r��l��9�7���w|�w���/� �@x���%��_���Zǉ-�&�
�%X�ߌ��c��L�87&6�
�������	��S�_�҈W:�,9�ڝ\)���X����I�z�Ь.�+�aŒ�5��h	V+ N��<��f��ߒ�6���[��V�N1�
�{��{
�����/�b�-�jf�~z�DVN3٪�H�6g,�a��>�]{-��gC^f<N�����S��;���N�"܃���馂�1�j�� �4�2�����_����T���%���|��}]��w��$f�[Cs��L-�bH���L��<uH���V�陕����.q�Dc����J��������YW[�P�Lٖ"UcN�0����:8Y�,���>���1[�m'��A�ӄg��br6k��%���],_\�4r��Y�%�=�43���2���46ǲ*q/�l�]����5��R�[�V/�R��W������r�ŰS��o��o]�����I?��?\xa�1�ŐUƳU�bUVf��U0ӿ�gfg���h|�i���|ҩ���4�~�o6_`��?�c�E����T_�H�p��2كP�Cd5����IK�	w�&�U�LIEn��[H���*c*�"wB�me+`���"�o��-�up�8 ��1�82��v-A,q��\�Y�ĲL'g�s��6��������.�H?��фǋ�f��7tܙF�~bfn��d����0�Y��!���;���<�aú�}jv���G�c�
	�:u�2����h8Hub�m�D)����W =�������:�M���`��q ̼c��=��J��
^bG�p�ω�H���ѩ�d>8(qo�A�b�2�#�������.'1 JL���^J_*�T$�1/ $�wӎ�C�')�/zыJb�;�����A��?��%�.k#wJ�F�$y�e��4���
���uի�l�N7�k���ې2/�~��?�ap�}�H9F�Cy��%b�,�Ԁ�^�{qOl��<�E�҇T���9u� <�L
'Oˍy����J�i���������v��� ��FLа� jf�$8Ǒ����庿�+�R���ჸ�O��O���[��vq�����z#�=k�[�\�$%�8��.h�#j�y�o�v�c,`,���H����g^���{�W��������*��C�y��=x�&�3�����Ek£�ɂ�����;�� �GԼ�%/*�����Z�&i$�<��/G�9߬:���9נ���C?�C�Ꮉ> N�Q�Z:��ِ�ŝ!��N���mk.[꺳��1�u���lǭl�v�������5b�`�%m֬�e����峟���(ו�����k<C���!^��6��]<'\d�� z��~�l"�����R��*`4/'��Cb����2��|�;���w��h�hŖ�C�u���3�3���@�u>5��'��� �I��饈N���[�����ϭl�v
 ����D�*�H��IOHk䄶RR�ϠM��Jk4i	�Ȑ�/�!1��#ΝA�l�g�XM�ݖ*���}6� �����/��n�����aš6DF �2 �/�JĊB���x�;�F��I 2��r��gl��w�hq�9Y�5;~�6�񻹘}������s2�7-,���=ϩ��u0V�#�Fw�c�N�,c{�ql�VF�tv��oDQ��qj��o��ͺ�j�uq���V�������}��ssN��E���ķĮ`=
%�ό��1���=
#�FFP�E�"�5�%����e�V6iܿ޼�mo���tB8xV@چ�Ù�j��􆚜D�(������K��`K� br���D��u2����;�7�r��sq�kC���1�.|Zr��c�tp��ǖW>Y쟌2��>5�&��C#mr�U���fƙ�Mnt���Y�ܸ-ʼg�Iw�B-�*�?�����'�z-[���8 L�b�S#���kv�\������:�g�t�u����l����?��#�[���t�E�<^���v�蒇DtX��J��a�!�u�B�X~�Ŀ�:Y��8x�>G�mp���p�R&T`�3:�B��Ӟ����;�io��a���0���$˰
~��c�mM���m�̳�U�;�ᣵ��sX2���(�˦��+RR� 1�Nm��;� ����	��o\Ì��C8���N[@JCw�`6�u6-q�t��6�z]V���	��4_�� R�_~ZH�0���LM
����?��>�Bl(���S ����Ǧ��h���)a���$˪P�	�����:���83N���[��2�O���'_oi��ՒTD����C@�Vn�ASŇ��"���.�ck�Uy��L���n�P�V�����P*�����r���v�1�Yˡ���>�3�Մg�Cs�lO9��sf�������QhN��fϹ���P�P�"�/���Pǝ+:���,j��+�A2�G�2���Ƴ��L��(GԂ�ГRpR&H��jBjdy"OK��vK u�d��mm�Q����8�9�F�d��}�{�of���;��P����Q��,J��q���2����
��#k�Ǔnb�݇�Eg֌8�8�bjV�F�\�n���P	��Eٱ�������F�3w;�l�����d��YR�uPІ,2~����`�@����ȅ���\͊���̫�3��]��'����r�d;ٞ��Z�i�G��s"��a
 �Fm�
�^W�Ns.y�[�;��U���cbP��!���$~^Y�&�|s0T�o���&�/sV�ɲ�R3e9)�Ԩ����N�8�&#�	W�1�.��!��%s�����9x�^�PVQjA�'��馆�3�6k���\�j��EZɶ�|���C���%WK�'��ɬr���K��y�_���r���s|5�#�A)�2!���5	�i�;U����4��R�]�R����Vd�^����m��~��_��(��v�9��`������t*�J(Hy��k�����t�X�����8����U�:	�j�`�8��LS|&)��RMi����F@\)J�E_�E��=���_�Ņ�$�	���>j����ٟ-��'8�������O~�G�p�ܓh�/��/)�d�
R��>[�q<B��ù8���?�G��	M�Yu7�--s������\o��*�-����F�i�;����9��V>Xƨ�C.��'�*0�O.�����$~w^Y��o��4�\��t.�1��̂�h8��p�2����㽒FpM*'c/�(\\��<v���J�p\^���w�� +٠�����Xw�=I��ⳟ\��c�[�1�a����'~∖Hb�ԡ�������<�9��#��ׯ��M�茉��a;��՟g[{~M�&�+fy��A�\��+�ͳr�浪�k9)S���M����k��e˺{��K>0=��<���Ϡp&h�
��L���J�w�Iih=x�4�r˗�����i��} w��2�vff8���q��X0�S��Z�E��aI��ß�q±V1D��c䀴�kh���1�9|�3�9�IH�c�A�A8�>�$�#���	�F�
��!}*z:Jk�RNP�.O�D��l����7�Vk����.����t���'�"��QF� �9R[�~�����{r.&*�I~�~C��ⰽ1w�(ը�q���f1~<K�;mHf�UZA�*�Nz,��m����IL6��	{-�<B]�P}����w�w����k���; �FIIYƃ�gL*ڷ�]2��O��1α�c��ˤ���w����H^���s��+�z-k��p
I-�ּ�9��Ԁ{���y:EM(� �4��Pe�0ǺK,@�Y�ɑ< }ҳ:�QKKm<�ޘ������[�*9λ%��2%Cǵڙf~�������~D� ���G �L�1��G]&�p.�e��yܗ�\Is�9:c�ύ�ВJ�t�j�Y���3lS۳NF��͘�\(<&�U~�S>��o�����Z�����*� K�S����.��v$�Y��EI�Ey������('�geC��s�F�A��	S��4M����-	&���~�`�4�k��s�A���:�z�5�Z�C2��.p�v+o�5��0����ukǩ�K:˱!�����*�z?�,A�E��������V���Nj��LJ���'>m�u/:E�b�7��k�YtrH��>Y6z�2v@���1�N��N��V�:�x���H���Ni =�H��1	�|D+v��jY���I���#��W�hz� �O�x���x����xԴ��2�;O�Im��ԨS�κ"��L�3z^��˒��6+7_W�������]��T�VaIM���*'^Ƹ��k _��%.x���Ό�'�Ho��7������\�O�o���E&c�0�:���8��PA��M�8���G\�8�D��ƩV0��� �1�P���t�5��L���>w,q�z-��'��I��*�OC`�����9�)x^���B�b�j�� �v�SJ �tw�����HW�{�3��g���4�l:�\rK3۹�z��<�ݥ\�l����E����OG�ٸnM��>H�8���`�[x��ɚ�hi��t�|���ef��	�p���s��UrA��v�Zc�T����F�{���fD%q�$@L;F��3� �"'5�V�-����w���^ku��U+���T�L�������2P�E��L�zQ�컼�3�OGlƆƘN�|���ZWY^���w�s���B. 0sE�2��2��4~��Oȅ�~�����N��'�����4���v��ݹ���{��r�nI[p	"�2/d�<WhӌyA��QIM�I�LS����� Nэ/��//�������'b�d]��$�Ok�KG+���ns��}?�>ۛ6��t��-��9�)��Pg��� ��D�	��������` R�/�K�3XX�X�l3\K]��JC$հ�$�w%��ꐷ\ 385�4��G ^e�
����ч����>�<A���@j DRK��p����XJG~Xm��E:-)�ia��-L���_�y$�`������K<<�s�g|�{�S
�[�tM�B��^Q"�S?�So��N_��'`��F��]�\�cn�mG�Ō����W��> 7[6�������/~IE���ښ� ��S����~����J�4 ���w$L)����%��/���{��	�����e�y�M7��r~�Yo�B�/9Ư=�ؒ�-Z�@8If�ġ-�R�Z����'�������>�nU:��j-hS����[/�d�ߵT�.Gj��P"�Y���5��x�L�I*$��y���~~������!iiy���Tº9ʱ�!衇J��ׯ}�k��ء�q
�K�x����QI�^�E|��F�7(@`���������e
A���x9 ���Z�A��r�8�[z�\}����>�SK�#;k��`�g����|тY�ȼa%�;���=/%��r?�Nxӛ�TJ(�n�V'�|_�_P��k
�9��l�U��xܛ�A}Q:ig��r�פ�>��?=R�����se�E�J$��=�yw_ϡk��ng�^fA8��4VDS�v�n���gc@q-��o��� X�TIJ����N�MP^j�`���v|$�'�@�@=��Z�H�@
C�Pm��pN�ǉ�%&A��oy�[�_��_+������%��X+0�(o� ,�E$�0Wğ���^���<P��^h�(��/��pٸ���&P)�1�+l;��M�Ox�S� n�$�x����Լ4{=�>�`���K�����<���/��/��|ei|�C�(���ȁ�N,�!��9�~k;^�nǤCE�L���8�a�����2#�`zd��r� �9��^k�h����\׺��,@[�<��Lzhk7H90��Eӂ3�,=�5�Z��:�2�;�65b?CR�^E{(*�akc�:��������ƨפ}��Ѐ�!N�3�s��{���s?�s��@��uH�� �@�{�mso����ŌfЄ/>:b>oG�Q;�ﴺa�y��>��E����������ұc\�������.Z-ׁw��0s`���W�������������u�5��ۿ��vr=���`�I��1�-�Ef1_,�Y����>��`���W�H��m�sZ¸]ہ����:h�<��a]�WϺ}ķW���x�+
 1���hY*lO��0��p��HWq�5@��K���\����1T/��T��	|x��_]ޑ9��7�qI�!���! �Ջe���i_��_ۼ��/l~��~�Ȃ��8ݠ `����Y U�2$�y(����;�8R�����^�L�I��:��p��Bf�<�'�q����bGs�Q-�FD�G��]�h(�;����
Au�4�4)���q�#��'I�tZ^���[�����ɖ�v��mM��l�hLLV)��t\�Wڅ�-��q�il�[/9�����4]M7	��0�|q�*][��W���	���F�6���^#�?3��Hϫ�jA�q���ь��]7G9������?+`
}/�jz�g�*v�Y�g��B�s��SN���P�xVh���������£#J�·jF�U���"X��qGd ӎ����P�<y9h	���
�'Z N3~%�/��\n��},��8�J���&��`�rq��g�.u0�q�d�����m�3=�I2�����dMm���{�+�fT���ٛ8'�r1��9�%��@���1� J�/�̾7�\^�qa8b��9�~g�U.� �1�>�4���u�k���ƍ�"�	��������jhj��,U�r��bA �Rp��4��d�{�myN~�b�9y/���vHŅ�΀W��^�aT��Թ���xM����vԍ�7�O���%R�/��/����� �أ!;8r[mX�I�ՄՍ�	��c�p��ꒋ1"������t�����!W��˭M��צ]���`�M��}��L+A 6D-���5���9�����x߭�:���e"��$����XT�
C>��`� � ���k��q�5���Z�
�s�I4�S��sƏ�w��~'���m�F�M�彩m̽P��`�u���=$yӥ}�
��O@5�����5�p�C:�td���� ��f�Z9D�ݳ\�&܎ǋŌ������%yHwS��r���ꏨ�f�$�J&�/�@W��x���vN;�ḁϲI���X��$�L��<Y���Y,��4j\�;��_?��hP���$t~~��T�`5�w�����$Ƿ��/����C��U\k��wU0��r��ߌy�_p�������,�c|y�t�^ř �o�����Q�Q$�)���D'�ǻ�.���,�/?mCA�6b�ءu�����}M���IR�`,%��Y+�Q��X0b��3�ɚ𸃠Yߐ��t��/6��4�SK�������CK`��R�v��0� ?9^���gpX�����zQ�Y�<��\�.,.����`)�.L(�52`~+�#u��N4�c�Ɋ���N��ܼ��� �J�;d�QFZ�^��#�d��?F�V�L�b�G 7�%�@��e�C�N�x�Q8(@��M�1�y3yV ؈��`��}w?��:-���W9@ՄYDT�2cϮ��Ԁs2Oǅm.qjM�ǒ�WV��<���e��ڹw��X� �+�����?���\��\���fŦ�����^aޖ`������,׋��]����}D:M�m�6t��5li'ʖ���6ʶC(/(
�UyWw#G��DH����43J&3��Y.|�Id4����^�4�|R�D�Pj��9��h���-�R���f�$�2��:�8(�����k��۾� ��~�����A��$�+��
O:@]��R��`�-�
�]��7:||<�`O��0�:h`�Q��R�e���f���������+��e_�A���(��� `��P3�s>˼yM�;Y䆙���&j�f��r�:<՘�����r+�+iN�4?1�	äo��˘Գ�Z�*mڟ'��B�T��7p?(�l	��?s���� -�3︟<�ڦ�8�7b��!��I�x��Fn�u��E%CF�K^����n��2��cwIg�JMǩH&Xg�"�[Z(����h���2�#�N؆��E01>����_:\4R��d;��A`�[�<�,�#�*�*�i�I=����Ⱥ�C4��PB�<����|6_:�)�����M�IN���{k	l���Em���(c葤ҩ�<I�J�	�1;�8s���"B>ǌ�F�.U�5��\���u��h�@F:��D����9o{��ʻ���>����P2���]��<3eP�W�+��j�$�����g�3��L:�J�?��c�D>���IZp�fzVYi�?�>�-�
���IEh��j�?�L~�!<0Vd��42���nI@�M�G�Nq�����=�@�=C��`�� �3������6�e�7z+�#�8a<耡cے�I���* ��;rHUf(�	[����w3+O��s&���q�Xs���*�������KA�����N\'�$܋g{��87���L�������,�����b�3D��YT�Ѩw��j�b6g�l'��h<-�0�>*3��?��J�����Y� )�j����rMz=��㚬pi�	@\�e/{Y�Q�F��Ȭ�Հ3f�,�W���������P��uO8���(��*���'��i�M[�3DK&)�4<J8�ag�(>g��%�̶�?����1����jق0���6��|��*@�ʔJV��Y;ƨ�\�|דD����zы^TƸad +��Q7Դ��-Fy�y~�s2輇�6-m��E�� '!�p�>r����k�	�%��N��� �>�����q�16.�A�`ry)_F�$7����А�wr�v*�!�y�k��C�;���0��?�S?�ܜ03��(M��e�y��̠2�Î7
BK��� 1aP�`�Y�t[�\Y�	�L^�P1��΅$-!�M�C[�\��Q�I��r[$5W~瘴l��� 67x徆�ɍf0�OJ�N�� ~9eD�.��8� �o��on|��bU�) 	�5�_���F� ^p<ֳ�������Z���%X��y�p�����͞A6J[��R:����L2L�O��Oj^��7ׯ�h>��?[�4���1�P**�����dU�=�Ƥb�����\)%G�Y��%7�xa;T�G�k3���@����9"�nQ��J��7*e�W�ˊ��N�\�5!�Y�G�8,`�NS��K���[���%#�$�o�"B,�W �����sė.�A�2 :��GY�s��	#�1p�`1GTPL쑣U[�Ӥ�zj��=�q���|S���Y  MFYB����u���
j�0������%>ڭ��ƿ뻾���;���e��1�F��rQ����,���r����Fb����5
^i�̦VM\����LZ�����a���d�����B�JY��O�����q`����6��%f���T&~�`��>v�&�⬐�X.iBls�r�i@;�lp}�\[���5��jIj5���8�@|���[��!���B��5r����A�t^�Y.�~�w�c�t�E"ǔ\*���sF$�J{dd��ajZ�|f�7c׹�U�)I�<+`��=�,
�S�V����=`���������u�ٗ���<�=�G#ϑ{?*�M�j��0�'�xtu�����_X^�	~%�Z ���Fc�Γ��@ ��uY�seup
�TMm��1���s@� �^�Z��Y������iz���j�i�aj���).Vj�75b@�j_��4uP'sMMX�~�1�Y_�- ���7���R���&�dn� ��s,�;[j�9�� H�$����AQ@Q�XY2V�_��Hh	C89��uZMe�IV#�|� �r�(��םj�<�s-B]��rĵr6�0���q����9��a�R���RM/�h~���<�h������bL��#Y�So,�Aʳf���������4�\Y�h��O��2����߮�6��(i�;Y��u�����Tn�%��EMg����E��4߭6|�Z`~F)V�m�X�:��R3<����  cq��q�?"˛r� z.�)�����e>����DI�5����\��ID%'��8�����7,'�����gý��wJ��1*-Fx���蘗�U�ח��y�CX��[k%�yoF3t�	�3q%�B��.��8�Y����W�Q_��o}�[�g�z�;%�Y�p��Sǂ�W��;��;CE\��m�d�K�!�J}7�h����!���?�>�1Ъ���-�!x� ߂��K�iMI�S��T�b_e���r,> �հDnnmeqr^�%�|�'�����ź��^�X3�6钌D�8Dʄ��[�%�㴐O9k�q,�<���:�sg񌭷x�A�0Ϩ�F`@�oJO��j����L�B*�=������7��1x;Tt��̧C
s�!ӱ�(A�����6��3�:�ģQ�D�z1��a���d�Ϡ�SNX��n ��q�vЛ�o8��9�,p#�ʨ���q�p�[	w���Ο�{ Tm13��.J-1N�qo|-�`h-�1�8�9f� (f���%c-w~q����_����n��c�z�'	mF���_���/��k[a��q���A8,�:X�?�EF����+�˱�k�$�������x|I!j8�\yv&}��^�sZ��+�������%����-���m9a���@q�M' �j�)ʧ���}�<8�L���Pc�����Lj5�h�	C?p�Zj�m+�c	��Nt���'����ݿ+��$p��4�jpy�:
�I�ǹ"`"����%�u9�,6��kX�Q�Z�>���~��o��r]�b���vQYWV�(Ƴ���F2�X ����S9�����` �)��iY�FP\��Yݝ�c���ɝfہ�������`r,A@U^�%M$�a!�& vb��� ���}�W�t��ۮ��b'Y@�Z�f5�����t&X��N�೚�C��{9RO��Y0�w�&
?L*�+�i�,��:�>S�SMm/�8X:�̮�Tz ��,c�}7��3��g��vN�$�/Ǡ�RF�9XN闬֦��u,�mq�,��s/J�I�A*ù�iھc.��8�xN��N��y� �Ĺ.��nz��>IRz9��,a�������&�ф�����軓%#4L�*9?8q&�+sZ��[�X3��)�#ﵕ��U���p�Ϛ��@k�&�"�R���C�{�/%?�|5O�RƔuX�_��{�Np�P�E�c�C�;D�X�`O��Ys�1��o�[`F?����*`f�|i��'��nV����\VY'��(�ssQƣҿ�ч�H���uWb�b�fQ��j��R#1[��;�ZD������V.Oj�A����c�!�t@��zr��
��HM1��R4�����ȥ��G����s�i��ؤ�q�=�������1ƽ���:M8ۢ�<\���(�~�����*�Z��(e��C��ƹ�dg��]܆9�(N&$'nz�kn�E*M�Ui+�:�A�OXT-5��H�B�֨\p9�T����:,��@̤���\�	��Ka��
�z�9�D6�Y�T�ۈ	�I� ZgY;Bz�{?���=�(-��Ƽ��P����2��q�^����c�&�n��� ��C~M�;�6�E�9�
�#F�j@��A=8�<�֞��VҏwI���-��c�41iUHZ�u�0 9F�u,���Z�TcG�㽾��ݑ[N@�FEj�n��C�{fVYf�%���]8�gH��\f�'�h�7���n.�g�� ������p �5���w; #�N�Bm�d�4�2?�ZH=�:u+�'�8F�'1�>�`� ������4r�[6��u#�w��Aҁ��?������+_j"�[()?ñ�ְP�Mm^P`��z�e(NIH���+�
�Wq��%�h�+5�Kq̝Vj �H�U���� ��Ť�T3�����ñ`VyJsP�N���H�' KG���/^�n����yV�c� sg�?�O���cܬ�5��rH��2�<���&/�q(S��2ؑ?MFk��*,�`|�r"/f�3��EM��#��}�� �`��"߭�b�tC��sn����\�V.WrqK>���2��H�7����ke�ǆ�R֞6�غ���9��v�����@VU�y�ȵ������PM'��s�C�;<6kN��:���JXu�Eʺ{]�p2O��-屲�1w)�d]U3�6	q��r<mb&��5�g�{��I�d�a2�I�)�U�����L��&��ˑ$
?#q���n�Ԥj�Q�5ـ1a�+=���6���ƕ#��qh��,Uh�E�.˙����sezr��Ҏ�t̩A�I���6$�$	������Eh_\4W|�ս
����6�4�ɸ%A�d������ Ð%wp���.��z@Mذd��9 WZ��U$�]}X/}�KK}
��	��Q�p��ʽ�61UD�\���ǥ*0m>��NI��o���/��|�V�c�=L�ɰC��^S.?7�o&��l�1`�	7�x����W�$������L4��*O|����
�l�U�;�l�[��)�Ǜ�f+گގ�	1?2Hm��'Z����~�k���e�;�ȝ5���*�H֡ �~��8���F�P��1@d�7��:/���;e >��3�[R���D��hՀ�:��G>�4qd�L�����_��R���g����4,/kf : 3�ٍM]��/]h<��f�fX 2��u�S+'���h����P���O*{��5ݐ�+]��s�� �i$�kG�O.� 3���Ea���u�+;�ґ=d�x�[����/�r���^��ׅ�$Ȩ]��ec��z�q�wX��k��֯�t���B�!�@�?���`��SǍ��u�Xx��q9���t�w$����K�dD��R�H�wr�逳�+0�u��3N��05A�k�E���o*9�Z�!o\�qc��J�*m�~G��̴h��X���:�d|��D]bv�aAr/F�CF����h�:2"(�Z����Va��#(4�3�E���g6�IJ�~PЄ��O�ce-'|p���C��bC��i�Xn<�	���E�ç��{�!��f��"/(�MU#4ƕdg�׽���m���7ӎ�B����z�j�j_f��~x�x�+W�݌;���f��3lĸj+��+y�ޔmۣ!Grq��j<��I�k���A.F\ۺ���1���ܚP.Y�$(�=���M�w�x,��ϡ{T�=��I;��G�8�������~��e����sj��t3O~������Sk6�LcK�q�x�(�`��;�V�����U�Z.����)�j)��\��I~����!������&Ub�r_+�Y����(�jÙ�9��9��h�`T�Q'ֳ��;��-�OGts����ޛ ݚ������t��!	�$l@.*�6(� �BDEL0�������[7Cݾ7�R�U^��X
j;&�hd0� *�DTEiA���3|�������o�o�=������~N���;�w�g=���4G���p���zsn8F�W��k��?�K(A��X�Y7t�L�=��O.������d�������Jg�@�T0�w�wO�Uy���������'��Ex�x0��d���K�����;��5��N�����e�s���>��W�bȓ����U��f��z����1��l

Q��I��@�Ș�$NA��~-�35�ǲ�����4�=X��]=#��X5'4��Ve�-��1WT�E�u�Y��H55�� (��/(�A��>P4V�Vf��#���ۻ�����\���F��3�)�ڎ)��Iyű�#_��fO^�A�7���V��؊��1l�]+|{���]5ƶ�b7�J����]߮&�����
�-E��*B�΢H;��f��#`r�z���������A�n��Ğ���G
l����,���:LT�Z�(�ۋ
���},�a��� '�,���9�sk��	 *��6M���gx	d?���}'Ha4�Co|��LD��r��,T�"� "�GU�fi[�E� f������e�Ls���-���w����.|��r,fgϻl��EH^\ೡ8�Af .+; ��gb�a�j��;M��	��K_�Ҳ8P������9���;4@�Ƚ ����<es�v-^z�$̆vk��\3������U�yl��O�y11�r���b��J�<�iO+*�z���7�,��t������j����z�"J�ű����ѽ�6�s,�@#[S{�^i:��À�.��%���/��0�j+2L���l���,lT;N�=��)@E�u��h�`L'�0��Ƈ�Fd���J�4�\L���	M��/���b�ӱ�=,��o�!� *���Y#�%5q%��Gi�RXr����q�(#ҙ����؏��t�2�r�P��"�ǋE�?�ma�f�/��S����l�rL�*�jM�j��J-s�$�4c�b���Y���ۄWV����䳞�����|�����:|�Cz@>,� A���Z�0P_�Aa"S�=+X�V
M�"��U*�c��(Tā��3)���p���8�m�'kH�����Z1�d��DӪt��չ`m��D�h�n#L���X�H��qW%�}����2OL�}���Mۅ�f|ޮ1n�c�b0�>_ބ BK��.+�ȍ?%~��$���c��Sё����4K�\�	�Z���s�8�M^�M��z1�o��V�	��	p�����s\{�E�
�D���at�&M}B���Q��R�L�{j.�A8͟���*��h�����q��Ak뭀�:?U�VWNs+jB�����<���p���8�`x7yP���v�+�+���EG�h�߻�S��.�t`���p�����k��%ӯ��������ӎ�;s�3�4md�����N ��ԩQ,zv�B4Mc���d�h��plB�9ǋ��mn���ow[��s\��"�[�h���X���7���T��N��b�SV�ct�)ɂ��ղ��(@�����\,f9���{k�P�z~֙�3tK\�g���6^�;}'�d�ۜA�~�`l����9��W���1��M{��z���]d��L2���� �)~�l�y�D;	���Eă�UV$�icU�h��u؉X�AԬv"?����HWAC�M������P��`�9��Ύ[*Mz�8��w�h6�S����6���ȏt��#���R�K�㱪��&B��$�c�H��`Z�k|��O?�я)����G�3���w��	�V���y�4���`�$�D_��ѧL
����3�!U\7.�f�H���q�F��lc"�4�-
�����n
8�4NI�.���~��F,��\�}&����U`:O���D:�;�09�w���Y<�ߐ+h�FY]��-����b�����ћ#�M����Fsթ�J�/�ˆ�A8�0d�Y�B�blN<��AxX&:Bt�Ȥ�qH�
����Y��o,�@��6�;��`:�cJa�6VQ��ɐ����n�v���X�j�B�	��� ��Ƞ�2ݽ��6�K^P�.�BȀ���n�i�;K��RMN�h��Z�g�i�7:22I�K��+_���=�cxG�Y_8��y��w�}�k���'�3�k!;@�P�\h>�}Ӂσ�%��q�]�V��'���:��3g�96���7G��PV����0l�P�����I�]疓8�aVI2X�ϱf:����0
B��;�u��7xn�3z\���H!4�j[e���.s��Y�=��7��Z}��L��|��2���e�l�{��a,�w�Z�?*���U�y-2��^���ٽ��,��DE���U���dY�}���s�}mҪ���~�g�h�|���F�#7�]6?�!@��_�C�r��aH��A �!�-��R�4|-ې�ؤ�L�0��(/�ى�2�'�^���5��/W#+si۲��0P������k�f�'I���Y:��/��0�����ogz�3����"���6�Ӆ	�&�&�D���03Q�N(��wm˽u>�6@������~� Nހ@�?�3?S�Ђ��L�:��� d@��K��<^I�\����F�K?DF������4e���]3ID��?����<��uו�c�E>`�@&������a��)� M���KS��nD���1��ʨ�9*�\Ͷ7�J�'�c*U ;6���������]>���-���(��,�j��ʢ#�Wņs�_���j$�E�μk؍�&�"X����*���1��ܓ�g˶�*}�_�2��q;w�t2�L7�dL��ݰ*�h[�\���X5��`a4"���P��K]LˮwP��E���F�(�(�^��-� ���_��.�i��o~sɠ���^f�M��Yo�vQ��v��?�M~��ʶQ�	�-�0�o��n���ډ�����X��)ҭ�R�@Ⱥ��!%; ��9�/� ����-E���5(;���=(�=���U�h��L0��Ô|�Ȕ夽h�_� ��hpb����#4��H��Ʋ�4Ҍ�=��@''<���U ��(���p=
azR�e�C��W���{��	c�	�z���9 ���E-�23
�N����N��R}+�Vy?*e���y,�	��[y�o4��&̱A<��
z�賙v~�'ծ���F{M�W.O{&�p����;G��_򒗔�#I���
��J�o4��{��.�S3��(�8N���R��a9��ن����k%�l<����`�C��횒2���?H�4�X-0���B�������B蘧V�� ��\�UuI8�įx�+J�Z��܃,6��sMl�fM��g�d��R�T���e��<�����i��-�뭴S��s��h0NW�;n�� .T_���<NQZ�M%�	������d����
c�;�!���U��&ev��?���k�gr�D<���7���\���f����na�<�ϻ�գ�������6����A<&� �Ǥ�Y�E�E6�Y8�M�����"G5fA���Y&�M�RF�)�c��(:�ع��}�|o�">�o� ������S�f�c�MԨ�>��h��r��-S0�{���)LxV�k����*�u�ݍ�zt �T��P�l�"4B�����<k��,B8kxʼzD�CN�ݝ׻ݽL�2���T���.�%]qFB�餃���R�jgdڻ�}����{������S%�����{
�#�����׷��嶟7'����v���+��~�n���"�����#$U�4���Ѱ���D���0���|�)�L�wz�H��KAݠ �j��5@q��F3�<�U��V������=�3�B��I&�B4lL���BK��6i �}S��i�0s�e>����~�b�G�^Ď�G,�� 1�Fަ��o�����^]�e��n��]�J�C�)@e����O��v�Q��ʫGgPro+�$�ێ��(�S�;.��i��e-{��8�����O�Y��/�՞k��2�D3��&v����,��A���pVPf�}��ש�h��qg��eV�jw�I!��f�x�W:��\h��wF,��E�y�����6��5�<��ܡ���%h�nLR��c�U#\���>��	��w�q�c�&�c*g��>Xm����J�i�I;��"4���ͫKt�g>�?�9�
ܜ��e`�D0�v>����ʕ��_��W��=n��꫋�x\Rs�tG�F��%]W�㤌M���z@��5�J�c�C�6��s�E�{Ht��̅ӱ��@�z�T��m�ud��, q^���] 8�{��ģ�a������ݑ]8D��v��6-+#ۅ����e/+�e����E%���!J���[M���S��a�G�Z���1�����\��SI�Y��-����	S�b�5��}a�6Cm�G=��%n���G�:�!�>(�/B�L94ˊ�	"���H���/.i�=&>uEA�T�'F�X�D����b��B���b��R���ksE�zҧ��ʦ��k�v^�7mf��QL��;�%师L�]O&�1� [�Y���A|�pD�����^�c�
�y�!� ��Q(���zU�D�Tl$s��0)�.L��Fq��F1�,N$?�W���V�>چ�=���1�R$��}��G�?�%������kvw� te�\�3Ep"����q�dh��"�R�[��L
%�9�)��r�������X�7��=>򑏔�,jU���U�z���/�ʖH�Kq���:k.B�ƐH �U��y��[� ��S�{��Jb-�=f��� $*��|Ϝ�t���"!� cY+�ۨ@��A|F���r<s�v�2]��y�5��(ؤ����,��M�Bc��_����D*f�c���e)Y�� %� SBa�[@����枤]�<�?�pݤc��6Gee�N��-%yb�D��続�?���.� 0B�,��at����A ����P'&�c�Q\����F3MWۙ�<M![hCU]�]�N�z��C0k�f5�bW���/m}�������B)l�SC����S�0�R�[)��ַ���[��"8���7�s$Z���b^q-�^��W4��?���LJ-�Ë\��o�!��;���M<>�������Y�/��/ԙ6�����ۿ�|�h �gĉfv-u"xVk##{�~]�X����h���g���ݐNw�D�`�@�q|ڝ��I+���Bx@�Q���&�s�O�6��qkY]>��/��-x8:,��
F��3�nR�v�D��M���6��Yp�O�QR�J�!C_L�>���ժ��n.�.�D����t%W}��R�Hdz�k��R�?�)�cjB9���5���(��Nt��f�|��8�����qJY��y��h�F"���\�hv@����|���)�!�)"Rw�ܛ>@���2������E�z�օ����	��Dv�!�耢s#T�5`���?C�l�Q��R	E�ⲫRЮ(%�u��Xcu����&HT%��4�cݞ����!H�ņ�I��G��o��b��ZT]���<P�5�3U9=��t|����"��v^��MӁ�c��^���)8�n��v>� S-t�o���`3��cR�}
��Qȝ!8�H�x�32�4��_CHQ�-t�-���)�W�)�ۍJ��`����h�����o�뻾��0i�*h8ܨ��%s��ұ�9}�s#G �`)���	�J<2�_���Q.����uD.��)��;�wW��JO�����>����ǉ��|i0O�J���5�#��]��0��~闦�`Z0^���A]�� ~ғ�����e�����#�fy�Y�e����<���y�9�	y�Ь~��T��\����'��K�~J6��o,��Ŝ�0��O����
#��bYF�ٽ�mo+�F��s 4�!,�� &:	r;M�鼭�$�W����q�")ʠt"" _f�������E����W�(R(sM^,PԞ�gʫ4:N.��$q�M�m;�:4LIU��ϕ���;褁�(��Ƴ	��0M���5�3�-��=�N�qڮ.��㦋�?���q��(h��;�EW"*�~���A�|��v;,�55ZH�� "~V�[{49��
A�����s�"D�%�a�-��=�g��X� j�̡4�%R�G
մ'_u1��1���_�j�T?P�	j�g�.���!Wڬ��a���bǪf�}t_�e������A����Ԁ&6e&�d���:�B4�ݗ��<Um���&�r5)�Paw��8�.K�b�l%�ˍ&2�Ӆ#�\��ϟ}��jW�h\J�w�!j[$ktk����O��X�+�fP��v��-��l��KA C��^��-37,b�KI_L��]�W��2�%��Ō�v�d�vv��������B=A���v�"h� �xf[iFМ��]��,@�%§>gdM�}ҡ��X�tGw�#g��hj0�]5��l��kj�I�Ţ�1��y�����h�B�`8�ť,����K���N쬧��s"c`u��(��03���:�����/�1<NT�����~�4�t5W%�ۧ�}�E�9zs���7��|)�0i����Jngb�_���6���Rt�]�4ϔ��|'�~���(��b/���rG���6�4a�Ӟ�'�iF�(�t �����^�"��xv���6k�'�%Q���ފ��޽9��"�Xf)�NR��;�	���g�-�� ]�,5̀�&��6;S�+�)�y�ܺ��i���,9�ߏ�v���*�j&�E[�_��[�id�k
_��)��T�S0�7?�"\�s4�n����s��m�o�t%"�p"Z�1�t%��e�>Ʌ� ��h�Vi�Җ���b�j�U#�e���J���,�(9���P�}��"T���lQ�z��E��������4�=}�������v�&2�kߏ)[��L6��!��<��|�WVS�f�-Qs��t�mH�q�/�ڶ3^W3�Ϻh�̣4�@�5_��OZ,�WT)n��q�6�>&�?*�i< �_j�[���ߙ5��VЋ��൬qꠤ�@�D4mx/�;Zd��g��8��g��Y���^S�Y?�(��e�Mڹ4٤-�g�g��يI�?���z��皕U���lm����W����LP�p,�{�>����e։��&e[D0�(������E��ϑ߉^�l��\�����Tצ��Od%�QH;o�
��i�NԘť<5/�R0j�����z{�4Zx=3�fQ �u|'�)��I>���=����{Q~���_.^8#{T���vA�H�[��Wzڋ�9e��B�n�p��z�R
�X(���T-j�!c�ex�� ��n�ݐ�\]�1�M2�� ��|�'���>��ƿm�!��iCS�7�s��u?���S8���A�/��E�6u2ʇ�s�ZX���m�hš���W�Q�G5n���J��r��v{啋���>S�]���9n�	B���N2R��%:�{��˩ۚ�L�C�Q^�k������	`��5���;���9g�f���U)s��Hj��>9��h08}�Hx8,����7L����[ؘ�v�^Yo��<;����J�ꖅ�U?\��xu:"�.Ls�/��m��-J�W`��9	jЫ<��|�(�A��\��������&k�f��j��j�,sRM�A��XMl+��^iphǃ�����N����ś����]^@�����~l,P��]�{������X�
9�,�(���@�xU���Җ��+?�b��Zjx)�Ҷ�ɝB@��e&��Ț���r#%��!�Ŧ(�y��ㇿ/���K�M��a)ۂ�^q�Q�#VVze��7��;U���W}�_o�k;��&ج�.i���$ۇL��C.0,F��6��w�@�E��*`S��d*�tl'����v�ʩ��DE
�p�B@�L�oE6�(�>�������!(0 �ͧ��\�Y⹇��t۰�V~����?�R�����0��֊ݝ�V����F�=��U� �[�M�sͥL���!��妗YQ�1��4�ɳ�δv�e�	XD5*�-j�^���IJ��m�Z�M>��q0o���0m�|��q�k�igتQ�>���"?i����]r	\S�%t����n��6���\!|������ŧ�����`�ln��'ڎm;���}�U͉S��yV��<�9�f�<t.e�O�5m�LΧCefW>�w����&�H�"�v���
X3�,b�03���J�n�"�SX/r�uۇ��b���R�+>��`d�Y2Q����.D�`/��������+��x��;K��,��u��w��޻]�A���ܫ���-2�a�p��=�����j+�vn�N4���#�B�����Љ>3�_��9���=c��
�=��%: �(�+�T@��m���C~OM��E�lw�-��kB���q�N�癙�TP�w�#Jfo��������������<��>�*(mY�X0�w��m�7ƍl��6�Q�_��<�1k�[t<<� _8Q�	a����.#(`�,jz�K�j߻�xgb�U��	��YE�Gu&��QϘB*2}
&'N2,��
��#���
T�B�.
]�*��Q��1��S��~�{��ez��B.l/%R�kʊ�ET���b۝h1�Z}p~��Э�쵼�}��f�s�����M�$x~����Ѣ�m&H�]p7N5�'O7ۣ����[��k>��ϵ���| \��=6��x��V���Xi�<��$66P�q�P"N����3�{�
�ź��l��`'�� IW�RX�9���k��e��A�Tf��o���ϥ�'���Ԗ��0s��6��ŏc�1���񿌜?��~��T�a�i�>��n��{p�w~k\�z��fY�9|�ӓݖ�'.�6P��qX���2��}m)pMiL�����z���m�D�aJ��d*���믟�.�`��&U�e�d:J���aS4��ך�]a;&&��|��3,C�&�'��?���/E�a������l�����Ye>� �F�w�£��o�Fi�y�9gx��XG��h�;c4ǳ=�Y�5�}̣���<Ӝ���f������|��vY�G���k����<�-��ۅ���͕ts~�b���{��8�΢a�x��#�wߗ��Z��@�0ο����h��O�Q����UĘ����}�X5����$+d���2������ȗ*f�����t�97�'�!��[��N�;0��^(��s�1��1�L~��~m��5�����/x��_��_�.|o��Tx��	��w(�A.���XC���:����$�7 �Iz�t�R�m���fj��n��mM����*���vyQ���(�/�R��~��`wh�ߩJa:����#�!9��� 08���9�( �+Ì8a�hv೓���A@�L��炥���h#��>����	R�fҊ��x�ϳe�	߻ןU��M��`� Y_�Ew�B�h�h�qeԎI�]�Ϸm�Ex�9��;����~�X�&�/-/��yT�4W�n5""�'�����>����~\�ܱ}�U�K�PD?#���'~�B9�w���uP��)���.�C�]6~jc���F�}���@Q�����f��1i�E�r'�e��|�3�Yd�;����ۿ���w�/�����R_�
6�Q��� y�<�AQ�S��]�R�����q-�sG�]I��+��3�	l������U$��oM
2��ЎRhhc���F�S:�� ��R�w����=�!�(�e�e��e�P�Iv%��%�禭++Q�7���P6h�E��̕i�Y�U��Z��2��6hW��z�3�'×�3ĉ��]sU���'�5�|Xkm[��^iE�U����볛줟v������jy�-kZ����Ҿ�a1b<W[�^8-�w`E�h��t>��4U�4�i6s.��N��hU��ڝN;�N!�b������W'sn�OĶ��&�;��ֺ���3"@���}��1���d$��Hǝ���h~q~z_��fJ�6#Tv��H�3��#O[n[�>̰���ꇚ��E��Uk̼�J� )&2���k�����!|Q�0=`�0�	"�2���_�I��P�.yL�<2�q�m��O鑌b�8�hXz�N����.���ҟ8i'כ>߰��J�ƈ05�o���$��L�a	^[��V���7�9�(o��֬�֊ѡ]^�Ai'�N�R�BL���s����"�ü�ͻw��-z�}7���X?�A��&�Ź�%��g47�tS�� &���1̽Պ]8�؇i��|�L��ҾX����eqWO6����9���
��z�)�^�$�r���s��PG� _lS\��VɬF%Cw1�/��y�<k����x�.�K{�I��Ьg�eJ�O
�����c43�tǉ�@Л��p,C�G�yI�W���N�a˞8��Rk�j��o����kMo@��N9��|�R
�Y<Q/�)h��Z�5�ݳ�"_��˜�ۜ'���e���_��c��� bh��ԴhLp�y�F���%K�*�5A�#�Y=��w@���	�ֶi騿���J8��r����)��N�C�U���i��A�a�����a�bl�f�m������l���`L�搮����Yh �LM�PD����:��eֽ�����i���f֯{df9h��[e��qZ��>�Zi�ޤ��j:����M����iX5ū5u�y쬿��,�t��� ��E/zQ�z	���# eK���ۈ�S����V�7��SKT �N��W����	���m��6ڝ�{mD�x�4U/8�g���C��ԙ75z� ^�4�{U�/�t�0�N�����jd�Up�Z�}���,4=��௙d����H��5tI�x��X}�.ҽ&�����V�)O�����D�p��¼ԗh�3�r~����y��^�ۼEt���K�*H�-5�8�)�&M	_�5_Ӽ��/-�  b^D��	�_����#������n��פ?'�(iZ��Fo�=�Ӗ{��c����	��1.�	Qgޘ.;�Q����ˈ�!�9Z����f����P�e4O��b�Y���N�E(��e�E��^`�۾���wfo�%�gԢ��T�����7,/2��ʫ!ss�����lM�d�]d��Z4��T�zQ��w�~�Z�C�JS�֏��-�B����w��(ur��~���9S��h�ܹP�����g��&�ű<L�+�}���s7����(-3�߆�X�^��f���?�8�D�؀�|��ߘ#>��UE�'g�X������y��"J�j}�A�<�;o�^��R#�"�g&�C��{�S�ؤ05[n����1KfX�p�����^��V����������fH�ۨ���K�,1�O�� ϲ)׿մ/Mf����z�����"��:l�K�/1�8�	�\��FL�<�D��g����6�/J�Ub��Od�>ZieоW��!j[#�sDz�w� �{P���}u���N�'RP�@)<�	OxBY�f�5�H�
Z,Ę��؂Q-�jA�`�+���v�SK����M��,;aݧyݬv������f\%m�B[��vnvz�6��IXk��m��ˠ�v|G؁����Aqᵂ�x��乊�btI��y�z�f�f�2�s�WW�ټs�^��j��"g�aH�W�V�ٝ�цMK�j��Y�7?ב^�-A_��P;X_/��hF��[��k�hgP�K]����n��������N�ґ����<xE?�яN�T���h��l v�uQY�}��t�����p��k���.2o� �>�'>��0YM���MR=i�Y��@0"ǳ �����$b��}�q��CaWs��ZG۹^��ELX&NТ崇�w���������4=ܭ3������I2�,�h֦��JU��n=��K������,B����nF�ԞX/μ��|s)Q-h�����^�ѵ�^;�D˰Ay��C�E����HL�ٝ!�y�i�R ��[��LQ�ݐ�=$V�v��;"H�'Z(�Ȑ��t�{lF8��7��M���}�ו�A��[��ɟ��TF�j�L�x5S�
]�ߝ�Y���`YQmy5ҬA��"��m_���<ٮ<��q��k�d3ȇ�F�j���|utD��f�H��2��!� S:�2�54�/"S�3�;�b�
�4�X��A�ٸ�����r-�d�Qf%���j2EڊP�Ǆ�/h/��xle,Rz�y7>۾6������2,}ɤ�=��Q]����λJ�Й��������R:mP��JɐM"ن�D1F�8���x` o�dʵ-/�E>W�n?���<ِ�����U^Ÿ�Y���"���k����M�y�{
����y��)r2[sY�h�\��0��3��̴�+�%1�+��υެIgh����xf��E�u�����2��H) $m�ޟ��N]ն_HЗ�X����3( �e�����j�S@%��]]�(+�)���+2��+M>H2]�\|�������䋿��(G�xP(�Zv���(p���I]�9 ��5r G+�Y�r7[&�s����X��s]�|��y�4���l{d�=���n}�G��eә�w˜.E��Z�{w��8q� tn�m��z���N��7�����Qn�4��(�jd�����V��O�������wi��t�V�V�B���|+�g55���u(HL1���� \��1V�Ԅh�*yV��!�3Y["͌������z�)/إb	��h��}�@�� ���y�\uQ}�D��!�.�q�K�Ej3i2��)��W�H�5���T@)� �m�D�(�G[M����N��_��_++*�"H� k�9�yN�Mj���R͟g���Y����Ⓕ�tY�&pPUwl{�^�k��.��R�rR��<�h��dz�5�p���_�+�n=�]���¤��2<�2�^,'Ka����8�����]dW6�;eLh\Vxe|͉íe�r�������M�Hr�X�9��7x������-:͚�FiG�R4�9e��B�ڿ��碑%S}>�Mm�9#R��ѥ�ڛ���"�5�P��ڃ %�־2?WP.H�P�P�Unh�Ȩ�Lh�����G���##��X��j�LS�A�DW�0�Z��&U�\� V>�T���&��*`�O��OM;S��E g�@D���m��Y��L&�h�{�*��".�q�r��$�x�h)LHg��c�J�QSH:I�N.�9�]h{��Y��[��!@���9�i���}�k]�jd|pE��q���cĿ3�)��z�_x�QmW;�+�Π�#��X�{���1�P�k֡�"��p�:s̶["��t5{h*��꼁rA�9D�]���	��^����������� P[��L���vhb��n��g�1���[�ȹ�};�~�GG,�'�������1v���f��Pm�H�,�a�h��a����ud�h��1g�2I��b���� ��i���\]s���Y�G���+�ղ�}:gr��{:F]XH(H�
�<�����a_om�0���ń��.D�����N�s4A�͸�Ψ��Y)���NwS.qÍN`�ž��#�7�C$/U��1�Ij�R�Q�m*D)e��X���s�\�e���^���ҧ /��9�����b߅�g�,�Bʸr�����e1b�	J��T#��o�ʚ	�j9������ZDN�;�>M��Gp��ϊs枳�����!'u2\��$(䤭O(��iO{ZA��z���+��+eP�v�����"��,]�=;�P��D�P)�Dz����<GT�0�ڳ��(;M	N��;�6gU,��ue�e��_
���{��p~���Z|�GeM�h�����[�IGc�:�.�}څ}�Ef��˽
���/e�ܔ��r�M;����B�6��p�N�.�s-CN�Ye{�.��{��N�E�<��gKg|���[%��p��/������r�Y���H$#"DЖ��<��!yuTJ��4�j���R�M�x�����4L롧�*Q�<���D߭˩
��4C;\]DPt\����o
9��5�)�'���Q,ЬP��j��^D�z��hK�p4�v-��
�I�v��L�k���Q;B��H���P��
�,l�ئF�t�jt�n�����-���&��m���λ2�<2�t��h��>z&5��?�-�A���d�	�V�����p�Slė2�����^�M>5N�hj��0�\�S8v	QH�r>A�O��(��U(�춋߻ڂ%����8��TL�:|F;��>�k��v>EE�ڴ���9� ��s��B�y��_�d����V%Ul/͸�֢sk��O5�U<U�o{�ۊ�Fx;6=�ڗ��t��b��	�����g���:���~I���T��ez�#QWmk��� �h�n�����=�jh��`l<�d�L�kT�.x�q�[���k������@a-�^�p8�y��F��C�u,뱆R t
�м�R�L�ؕ�=�G�]>��8�H�D��x�͋_���)OyJq�s?�I�"��L:�dSon���<LԿ������s�S[8u@�fd����P"Vn�=�F����Fꕖ�~��)�)[���
_h?��yt���4N�m���w&;p7:�,ҥ,όZ����[�����y Ӽ���E�%�XcзU��ַ�=X���B@S_BP!�U�.k�祶�5 ��4y֣������R�ⶻok>��6w������Ul>�'٬�Ϫ�:�h�����I5�T�ۢ�v9��J��$����E�y�7)��w���σ}�t5J�t�u����O� �2���1�"{��V�yx�m�]4��}i��j�Ӷ�誨IS'*�*1�S(���^�2J�b~.��Y��B\M��y�Zi��4£�e��Y����2�Nc��[�~6��vK�ܼ�&�M��_p�K�q9�aA�<��z]A�~�|
[Mځ1I�����S����e�i�ά`���#��hsí�R�l�����D8����T���p�ݦ�Xt��6v�N �ź���ric,���܅�b�OA�^�+��f�ʌ���[o4�s�pυ�.�t,�5^|-q�r��dw�@�Z���!�4h##������y������<� ϸ���7*��iW��v��}���-��<��YIw��������OpW�e�?,]�4)�>�É����5��񽴷�����l�w����d��y�(��D���0��Q[v���0��cȘk��m���a��/'�?Zj�Xf�Q���X?Lx0KlV��A���Mx4)��Oa8�3�F��E,8�i�o���qͯ��U�ƌU��+
�Ġ�@9bA۠��ݬ���e�_:�2���zj�I��7��w���dS�f����]F��r�ڬ�+�n�E+Ee�V]Z�;�����-ȳ��kHa�M9ߧ��Aa|�tX��7��㘳��ڂ35�cY��ΰ>� �L��GQ�0��u�	K�LQ�暃N��)�ks��ze:m쾬��ԟ\�ܹ#�,cc?!��(6b=ތ	������'��~�p����3��#��a�'�2S���2� ʪ���'�����[D�c�"[^#�-b5��a͸�	#�<��7M8˦��	SE�Wb�.�8 ����/~�#�����N�$�R�	 �;�9䠂q�����A:
JA��m��2�明<K�@"E�נ�eg�Y�59�FK�#.'��z��)#Q"�6�E��2�3ge���A��I�>�@��d�Q��F³4;�`���s�w\����1��e:�h� �}�0�=Z
s�tJ֛H�|�s҃t_P��*!@��=�n�iɐZ��Y��g8��i�.{!��D�ڈ�,6ߥԤY8�����R����Z$�����dĒ����^��xt�s�q9�"a8�zT�.C�VĂ��fM��`�ti�|�++�e�4=d�nskqw��A��Lz����.{$�l�3��(���YK�e�N]�X�=��=H� ��-k��)3T�4�oC�F mpt��� �G���W����]֮XF2��8m�҃t�R]WSD�,�G��eM�4A̪i�`��^��0dQlw� �(�y�Ö���j5~�#�K��N�3�򸖉%x��u7ǝw
O�@O��-�Q1�1�n��*b�Z�Z,��?큦�&:�Tt%vͦ&+�s���O�B�X���7E��	kvXa�ο�[.����g=�\볟�ly���}��ԧ�xn§���չ��Zͼ~��G���_��e�6�~��X�Q'+�j}A����ig��ǔ�F�pj���Ju2�	[1�0�e]����u���S@]A�߅��~���wwW�L�L��N��v��`K��
���3
����������˱0E���暹����~��C�^L�����^َ�Ҝ#c~��/��	QGR�H���]OO'�&]����~i/�X��)�ԏ|�#�lN8ⴟ���6Ox���}�c�w~s�F������2&��{�W���r_V6d�~�~�,z*�]�X�RO��E���GuD@�-vM4�Lهf�AY;���4#~��`,��a����yO���l/�.6|����y�K_zA�^H��w��쀮V�M��Me�,��q�-6�u�u��L1���C<:�I��")�f 	1��l�����&�Գ�W�Y<\�Gx���!L�!��gU~h�������w�5KU��qYr�@(���-8��)w�6�ߝ�3��c���*Z���,��g��1���?��JSR]�oY�.�ܭ7�??/"3��_7��><�a�5��nj����<7�����٘<�n-��b��\lsOC��eȚg���u��a�������i�^���ovmI�0*C��=���뻦��D�	  ��8��H$��=*r?����]�2!�dr��
=�e��d`�8N
�Da�f���@��x+jy}���+�Nn��/����_�����Yί$c�	'��.�ۏ��$"�V0��\Y�hrh�ews�r�pr��Yu�_}��g?{�N���N�c*J�T����+['���~�Y�A`$�U[��� wa�w�Ff�~��8��b�
(�͢e��V��q8�D��s?�Ð��>5:$N����~N��W�m�|ge=?���^J����C�9����sKV���r3�.�F"}�e�p����	z���wP�{�s]l�hkɷ���P�U�Ml���]��1���D�����`��,b���P�P��-����?��He����-������� ew
8(��JN�܄�3��}��Y^�.H���18�D��#%���z��D�j	)DT�sgm�:n�Fѹ�0��6z>�0�dͣY}4K��f�Ft	�d|<^j�ٮ�C~ss^(5�	G����l����D���D�:��oc��un^+�v��[d�耓���2�L�JS���c-]{g��9T�at��ǧ�`2!�q�bR}��xGE6��N[0�0�Cާ����� Ƴ�Șŏ������|���k�A�v�5�R��9�g�g�3������|ڥc��>�f���O���J��K� �3�Ф �G<��g����~y������s�|����s Pu��ϴ�g���s_Y�v�絉ľR�+�E��F�h�j�-��OԶ�h3��^��q|VD�����s��ۜ�v����{,�Q�1���p����&,RϫW\d΅�E^�d���;��LD*L}򓟜��yԤ�K`1�;����z�.!Z��mևN{���	C "PR��!Pm_��W�sElLZ"@wD8�������"-=����W
�T�^� �DB�ig�G��ɾ�Mܗ��?��?�jg�+�Ȫd�k�����;���R�3�#�+���s�M<�O��2%�c��3f�A�"���[�G�Q���f~�nL�ᗾ���f�����h�pck4?ad⛕f�4���V��±ߞ3��KkG�o��x߰��h&;4􇹡�{뎏N�=�sVBp�"Wk�뮛2h���e3�*C��V����t�pkC21�a��z]�r�Z������Y�&K:��	�E�$t�-�w��%��g�4!dZ���6B�2?��?X���C�6M�lV�cr���?��?l���7��G����YD�=�=9��p�'=�I�����s�."Q���o>m��2�|��6R�xj��4��~��ӟ���ܐX53B4q�9:�k^�{���d����VB��dK������*��3�)Z�&�vv�K�0G.t�~^u�aj�ӄݖmͧ;"��+�&4
�f�����q��^�"������+8e�D�V����Hr?<&2��C�MU��J��Q_;횵�Lov���I�9G�� v�/b|��V��ޞ��t��6����
=�^���1��z�0��8`���3M��D"8�ːp�gد�_;�Db����өC�E�w����ɟ,h�6s���H�tJf	J�r�]�j���U;K�gJ>�\�w�jG���(�:�Mb)Fnm3i\iZ�MEq+x�F�oƂ����u��|��R��C����=�Π�*���_U�z���j!�9�"a�y��;0�,A9w��x]�Ʋ{�Tx�|f�i�4�B��n���&��ϴ��c�� �ڎS����и��+
ә7c7�CS-���&���h$�h�UՇ�8���Y6��]��[��NmNgf�ʛ��ߜW��g	��P�	߳�9:�ϋ�!�	�~�}�N��p�}�!P��ឳ�!d��9�<���u2���
M�sʕhmV�LI�W�0��=o� �����<T� h@���f���:B2p��`QbrY�6�Q�i�L�,�I_�r{�e�i)HLڊ53d���g�`���r���§�6y�g�������l�;�<��7������ʃ5�p�#�򾦨�M�}.�5_�}s���t($� �Q��v��W�:���2Hw8����>lrw�r���� �������nj��,A��9�\���Q��ʛ%���.�!�������jXm���ѿ�g��o����x9l��`9���:�>�Ut��G�gݍ��{N��B�{�Y���i.��I;n�B�Tq_]��}�B�b��3u�^�1�Ye�� �\S;�o��1�����Jm�>��}p�f���N`ϟB.c����p�ĩ��#8���ۮX�G��_��E�m��0���Ɵ'N���:El�z��C�[�Wځ���������O�o6��@H�
(��#���^��gQ
�d�4C̚��T#s���F3��,L��U֪?����xS0�M�߬�����57�!f<�QR��]���&���|� �@�X0��(���-.�i�2t�"K���Zf�5������E?��,�̉y�y��xl�.:(�Nw���vk��lU�MlX��c���5�=(��{?�o�3�><�.`��x`,�/���åJW�g0�H�K�Q`��[����x�rY%+�O�i��N�ɬ����s-��~��2J4m4��`GmT@&�M�B�&�	�̊�j�p1�q��fۛ��\��!�+�k��7��}Ώ��E��������?��D�T�Jy���W6����y �v�)�3��1�:��@�_5�4�0�,X����J�����(�r9
�Y�9☣#���(Q��nc����u�f���$���Ex�&��oW-|j�ϴUVz�?��&4�I57S}s�s��~��e"�ݿ�w2�5g{2 >C�2LG�Fĵ��ZLG�舮j�D��h~�F������ʢ`C ���O�8y.���^N4eg��Z�ǋv��s�S�h?�<J�-��<��գ���?���������FG(|�9���Q���-K)�چY��5A�)B��gj��>Ke2�Dg ���K^��/3�Ĩi�)myQ'"lGC�	�"���U����F�������Yk%iq���-�poT�-�r���������=G�f|h���8�d�X`l^��;�SJ��=7=���f��ZAo�ۋ�&��	��-T�^�{Eo����/=�
*l�L�.{�#p� ߯��B2<�'|*�ʈ�&�Z������o.P��Ԝ�����e�b0N�������O���t�!h�P�i���<�'ٿ��d�x�[���t�ME b>��k�����k^���6�Z�֋�NJy�y@FZ�}����T�1��L�X(k�A�_�ѧ�7���T����˄�t@�2�|�䳎tqBԦBvT�cy���٪� �^�R0#����� �ڼ�v`OA1��>���
C:og06?�W�5~�}�v��?���bC����N�-�$�����P:�r¨T�m�p��۾��u�ٜ�F��o,�h�(�XC��y2����V$l�En�äE��2�H��C�d5�ְ*kB���>�<J3�Q�}`yO�^�	���-��@�@���f����@\s� �T匚�|4�v.�y�.�4M[9����7�&��O��V۝ʱ���s�����#�A �!ad�=Z-6�V5;�z�[� ��I������pТޖ����j����V���V�A�c#p�fפq]�`bׅ��i�Ө�=+M
�����h��*��I��@��G�o��h&���� kRNM@������M�]ǂ�W�����i��N2�j�Ь�DTƣZx��07�
c���|hz���}��i���f����]��a�ɲ8g�	G���?��X^�A���w|�\B�R�m�s��yF��3���:W������3�Z���w  ���,��u�ˌIx����#�mv�X���j��;=�\r�
���b�f�����l�����6����VVWoﭮ���6ۡ���������p������m��j��+��S뽕��5���i�;;��#�7 `�A2��	�l2���5&�G�T_p���*�I
��x�_}\�cQQ��X�t�+���ɿsҙ��9 :P��j�E�u�tMYD����O|b�7�aϹN^�Wۍk[�~��㢌 A00��ء�i|;�n���	������_�*~��#�_d��\� 7�P����r�"�f�X��v1R�b6�Y[3W����Dۘ��&5P�
f}]�އ�%��9��bѝ�H�`^�"��k�g��m�k'��ub����S:<q��m��S_X;ٿc��~��Be{pb�3ē����G�Νy����Sw67?�<zg�������U�Q���';E��q`Pj;Q�l)���t]A1KT����S���*t��,�嗿��͓����0|�[�ZTP.�T�W��_J��I&���,2�yf�!ϯ���'��֎Ό�p1L4g�jީ�6ե��%��Ї�Ї
o��u�+� t��c������O�g�9E�:K�G{Ws�}���'���?}"��'��yâN^��m���  G�\��d�A�ӋBY��P�m=6�����@x�I�Y���w������^�������m���W=䃽S��sW��~����}��Woͺ��7�w��ӟ�X���U���Ǐ���g�~v�̝�\��~�a�!�ع��g�_��Q�dK��yلt�#DE�:�p�Y4H{h�MoFmReco.���;<ݿ�˿\�b��>�,�js����p��F�^R��tX^"�e����?۔��*o�ڋ�~�2��~����0}I\�/��/�=E��vJ��K4~�߂��|�0��
Jx7��E�6��p�s���31Ͼ�[��h� b��)��
��=�s'�o��oO�AF�dx�qҡf1afTI�o��!����k[�'O~~p�C>�y�U�>����g7��I7��|F�י����������?_������o�>�՝�����>��1��Xg�G]�&�A�ƫ��1�9�����_}��W��`l����jm.�����8���>�,�(��o3Ѳ�/�2����p���z�긓>���x�R���ߘ�@r� �qcƯ��l���4f��� �g]5�״�BڬYl�M!���E�"�se֣ a����0��PW�Im��� ��"��	��`Yσ8�<Nx�<�茘Ҟ���<-C�O4�VV7�n���֕y��UyO�a���O���es@������z�?񾇝�����'���yp��ן}�7��5ɬ+�dҍ+�MPڴ�İ��F+Ӻ0�[Y��U���:����Jʤ�;���
�Y�9�<8XP�x�ɬ�ʻ�L8�u/�^���$����\}C��&�B���{�)��Vp���l�"{�bV`)���ؤ&/���3��50�]_d�K��e�R�y�o�PTô��8����!g�S�z�э�ŝPCR�+�^XD��1�e����>���2��S�G�	���˦�&G�.K��y���P[��h�����8��s��݃��������}��s����?�����So��/6���hV������+7��*4h���v5�W���_�����f=,��$ʢ�g�����ZA��ŋ1�:��Q��D�:��^&m$��«�C���6���Ѱ[!L�v�N��2R𤗹F���Y!j�'_���8��Ƣk{l�7Qp-��]��y����1HMH�X��6�d��BH�b%������)�B��O��O�1�
J'S�^)�f����q|�jkj3�A��f�5zh?!`�ۍ �������<K�]����C�e6`nQ ��^.�z�<c��9�6:"i4���������t�ݜ�m�������_y���C?��׿��8�������/~�CkW>���F�ίYkzW�{L�Qz;�����~��8Iz��W�cw���ʇ4ḁ��l'[����؛`2P,�N�y�BF#��UY'�s��ܢz"��&�\��
�+��d.��ȝlf��f	���RsrմL��2��3/{>��
%��k�~��R�ÏV���L����/�2 �dLX�+^���~�Ǧ��2痾���ق�O_�QD�=��y�5Ρ��,��c΢��B�9��w�wO��C.�5�����/�����i�maԻ��	���l������s-�:u⏆W�~���'��/nx���1�-?��}�i�����`�����\��5�vm�[/��j�;�bP�K,�����|Q�e�7n1L�BH�Gm�fM��h�+91����w�|�+���+���#g��.θ��L�]"��Х.d�Ѭ����P-������\HDU�%�	K�"��^\􋠂� 8ٺԾP�����7�\�ז�(��HQkk�ׄ�y���β��"a�-����x�k^S�jS�AHsJ�f@栵34��X���Q��Gl.���j�_Yk�������[}�G�u������1�����������7���w�����7�|F�>ͥCc9ܯ&�pƼZm;��xFab:�TH�1kJ��^W	[�{v6ÄX�l�|�:"s� ʁ	ͱ�`�~��KFcEO[�ahV�X~���c���}�s*���lbR�Ǽkxy��	� ��Ř�)a&~�@��)'��3Q">����j��BV�<@˃�A�%��>�N�����%�A�_���xz5D��i7f2i������훠�᱙#�Q��0Zoz�'ϵ�����?������>��+��k����:�I+۫덆'��z�qt�Q�+��F�J֞� �|�b	�1Y��v�%]�|9k������N�L`������L{��f��]:K4��%P갠K�RŮ�(tXD��<s-�<A���sSP��=Hm��P/Y����wY�s��� m2>�!�KPt�9�O�������p���f��F�)Q�O��@^KM�P66���_���1�>�~�0�ߏ��Go-�-�ڇ��F<�/����=�~ss��7���'����GW��9�[��~�~e�k�hX�hkL� յpxY=M䒔�c t�������EH'w�5��
��|
g�.*�Ӗ�m���1�����.aH�h��P����&lȖ5��:�vQ�)L��&<���}Qɩ����6�%@�
�.��������9>��@����m�s�B����z"�Ed��@ �`$�>,�98��>ۇ��h%�$�����տ�Վ��3X?�?6O�x�'������>��kk�>}�7�����`篍��2
+X�{��E{J��1q6YMlĮ=o+�&ֶ�M���%9X
\���SebtCdtr-�I2�L]�EyH��ѱ�%��`wCxX0x.P�QT����R���j�zm�?�Y%���+�.�c�V,ͺ�ـ���O�I�L� R����wO�]��귄���h��)�G�`d��،E�HF�:7Zլ���|��˽<f�7,2����}��U4e����Y�F�n����룍Sw�_����ɵ?k�c���_���'�|���A���͠z�'���kE��}�c�⢎i }� ����sY��\�A�;�
VO��vf�>�/�o�����ȝ!pȩ*v���\��Q�}XA</�������2+�������&������"�1%���a��ʐ.$D�5Gl�'�$�߬{��?&�5�a�8�ۺ
A`E3�&!��I�hl��qaX��25�,�!�b�@x��n;�����`XP01^�G��&t�q�c���� ������\u��'�z�؂��7���a}�����m��k�VUMV��N769�C$���K���-T���:Hǂ81�����b���$�)�c�Q�Ҹ��yWgse�a�ߨ�˖1u��lzk���IO�hٰ�>�$Fp{\?�2�5�@�'Nxۤ����!?NJ�������ctpZ�ŅqY���^��F0�k8�ue�H�X��E��'�s1,cK袻m��rA�]D����������_�k��5�3]Y7��a�f��7h@�]�ɺ�j���?������X�MVȲx"��{��8������Bxp�Lo��.�������k����$e��++��N�E��~oog��a�h0��������V ����1eƆ�X�(D�M[��ݔS-�z7[B�s3�;2�B��Y���jS���߳��]��\ՙ��q h�:�U;v5Na�=�+�<�XQ���gϻT���?�JAg�%��u��l4H��E�3^,���-��@ծJ;�����,���R܉�Y�0� )���h<n��ŋD�P:ʠ�B��VމYw�E���pXPh'Z  �hX���C�7{�:�4"�D� X���w�I����I��^�J�������-�l�ߺu����DgO��w�ε�{��{)]��:��	1��`�"��&Ӹ����)@a>L
xuq,�P��}3�����L�aT�5�!�,���.����H��:׈̐&"�ﮓ:��tI���sml�81��=�=��y�ѥ �]XV>+�8�9r1�8XȌ�YV���׾p6��q�Oe���-�9��|D'���G>򑢲c�!˫�[A�+���H[Ԋ�%����E��FD<^�f���C�-`Ig�<^��M���nIu�<����\�?4��W�7����^�k.�nN�������B�e�$S�����%h۽1v�3X�����3 Z<��Lm}���3S�r��tҩ���`�d���U�d����@�.��䟌Օ�k>�o*��%�f����T2�jDs)�Y�M�x��������3ĩZW`�"�w�g
/� 3�Q�[�����E`cG~ӛ�T�0�������8�>�M�k�4���j.�>�s��\҃y������C�����u�ڡ�f�����Ͳ��C�{2wj'�QDAkG���W�K��Ѯ��;m�Μ���x�7�AU
�*Lt�9b���d�����ΰ (�h���  �3�|��nGt�(��1�Đ�b��,�D�n�.Ѽ��i�E�h�캚�!9FX��\���\��k���)�J�J)�ٯ<��3jf���������N;���#2US��A��A�8;3B��R��{�w��r���cN^�9�ݐ4CE�.X.4���_�Q
�@�w�K{��q_�s�>H��:s�r�>����oIZB'}���]�Z��8o�oj�mtP^����6gϟk�7w��u��n���X�q!WhQ�L�<�o��Ewjǈ��w��3%�8��f��	nXS^6������4mc��ն��K���ڜD����J��մ��E��T�Q�=��nl�p��U��1�Y��EW��w^�WcsQ,�����k�(��.�FZ��h	(Ζ,Ma\/j�0�9#E���]n���U)����0�n%Ys�*0���67�5����Q��.vd�?�wv'�`�[K��Ɖ�ϱQgF(�\�Ex2�B��PX�nD�N�L<Q���N���zO/z�	���qMuZ�bׂ�5�3��U�\�ḿ�lӌq)�$jS�@��*3~T!�y�ť��86
�T�6@`q=�-�s!y����F�i�{-{�qHZ~Ja�(�d\\d2�85A�a�^�v�<94�qmHm�y�}LܨX�;}<s]��vv���/e�;� �V;�KK��8��Op)�n�C��B2İ�ӻ��n_��t�Wl�ﾲ]OW}��h��zŚ��u�9yb\����얦��k���6�O����Y�r�2�,y��X�tR>�Ne�I�3M��5�)@Rșƪ�
bJ��bemUX�>�̉���&����'�Œ1�
)��M6A�]�KCyF���(o�;�S�)L�\8���9j�>1d�J���|�}��rGp�s��!�O�N?F��8�|��WM=���!&��7�����"�;�`�~��߅�-��Rk�2I|hW��N�-K5�щ���ک՝��lJ!��}u�l�b��=o�����iVڱ�z��f�?.a9n7�_h�����y�U�ze���kǵ%B͑���~��D
�Q��r3BU.��W�WK:�ꠅ��頼_M5�f��~��|�Y�����ɘ0�uT<�H8mԗ2�N��3����i����C�{�!f)D�Eϩ~f�L��-o{�ۚ�����X򥱻����L��@�E�<pw�)of?)�r;yy-#0܆`f?��8=���:��ej�fa��h$�
ND�vk�Ȥ�Y�&ΏI�(uo9��N�ܐ1���՝�W�v6�����W}�E��}L�;mek�-nX'U�K_�vƥ�餭���1�	��i����|3l�J�vONd�	��L[����)%ӊ:-��w�I�'[U�+��Y"0e�E�:Lތ���)��>�L�^tE�])�:�uĀ�a3hG�8�$`{��ҟ�fι!���󬝒�D���~5H�l,zj^�gTK���"&�s׵�Y��t��4��?5O���Y�n۴�-+eN^��n�������9������P<���7޸2��?bo�����G�b8��XN�Tk�V+�W��ca<)�Xl`-���L�� �T�e�E6[3������L�a�rɕ�Fl���TSiY|kR�	�ʐ5ⵄ⥎��t�9!y��+��LB��/��4e9~VJ#L��<��$�m�1m����?���~�2�NH���z}ۇ�i�S"���t��Z�,���0��d�q�K��~����9�1�_γ@�7��	�T_�.�M���y�c�C��o϶�̭O��x�Sox�g�n��G��[n{�`�oX��z��p��S �v��={g0*q#'Z����l6'N��
K:[���n���&		&�� ��E,��'g�&�B�(�(��oJ�0Y��qN��6[���ښ��7(٢.��3.)���:4���������^"�4}1$< ��A#���Fiy����B�*�3�7#���1P�1�����W_����d�l�u�!A�fO���:�Ut-�ʵ��_}�u��a(�Qɳ9ޔpg�:V�(hA/�:n�Ȋc�z�L��k��Z���湝ǯ�{�3������o?��t�����k[i�5+��IWK{�������q����x[txr�9��hΞۜ&R����|`�	�gr�s�A|�63�3@���|O��QM�U�Yq���t���`ڃ���q�v����Xe.�
$���}�R%�!ǖ�s\ja�3[����a��?�X�чSM�EC�|='ۚ��4w�	2"Pڥ=^���w��S�UѪ܍E��-}������ c(�ǟ�n�s��/#���ģ^q�"vX�E,�cBA���KKZ�K��^��8�4�L���7��S����{�I��g����n�����ǭ=�Qͭ�]��u�	+Ý+Vʆ�Â�K�{ㆮ��0��j�`�!���:�ew��1��wu��g�&���2�67�p<dc��Y���r�6+����</�-���٢{��D���y�g���R� ү�ў�����1���@�2ce�~A�6\ZO�Y%b�����{ɧ.�6X��s���cjU9?D�"�j�P+�gN���A$��G�8�wT~�\��Txjrr���>�*j��'{�������Qq�x/K8�joxf��;�y����x{ȁ���D7޸r��_����OY�����!��m����R-Z��C���v�J��F���V�����g>5a�a����0�^��WM�����R.7�j9����ľT�&��ZV�ʭnCi�K��3�A�@��0���,�d�/��,��Җ�,��)��Dڼ3\K�flo��B�q *�%���X�y^�6�ϐ*��M���وP�
CFBh�b7g�0��n��E�Ĝ܇ҕ��sσI�~ꧦ��9A�u&�9/2[�=�m����<ƉyTk
a��}'ьs�����rG��h6Z9vb��Ki� ��Qg8h6Z49��z��]�|ss��w>����^ks�
�}⎧������{�z����ںN�I4�8ך���Ѷg�}��hՉ�v�yc!Dm����)�Rq�\}3��>�^�Bȩ��(Ԋ56��`&���ht�Π���&`V��v>m��q- D��/�lE��_L�h��?j;fF)ty�DN^���A���O��6�'��6��ΩN���H�
��d�M�cY(E�)K����v$1�!\��S ɬQ�T�KH�����nsDQ{�0�uY�uu)`�&�v1�0&V6tN��c�X�O�*��Ѱ���ޠ���������i;u�
�a����gn���S�������7��?>���Z|ݟ~�/����/����x����+(K�&��+po�LG���]��v��y�7壘�D6�3�©�����Pb5k��P*�#/��mͲ���|�̧J)��ȳRHUJ�q��j;�1�-C�,C�	��6�@��E����h��{�Yז��ꈊzLs��̞T���3�*I�1Ρ���uf��c��9W�N����]�]���z׻�Ü���ٮ\�R����	�r�1��t�M�(�u��i�����4j������[]+[����Q;N����͗��h�;9>l��۞������������w����O5G@W��3'N����in��[7��E�v�>����:��~ �����}�mF�gt�T��.�<�Χ?��� TO:�dl(F]T�ļ٤k���0��&`��L~��ɉ�3&��E$'oz��=���p.��E�BB�f9&GL,�:*C�xT&��M��qн��on^��וJr�%���X2Ь?�׹�V���o"<#�����|Ԙ��Z�?�ݖ{���aoeg�26�kK�o�� ���ŃV�g�;E4���#���z�+v��!?�Ʒ�x���=D��k~�M������o���7����ۛW���ۓ@�X�܈�"vx������͸��|�T��F�ZO��R@�z�]�ݵ���|f	���11E�:���oR��!Q�IJ��	�|�/��5�����늶1�Y�1��yη�LEN�./Q�6����}���0��~N�0��-oi��ۿ�b��pNa��w��1�sc>!��(J�v:��6y���< ���
��;->?�vJ��x�L2ϲ1�p����J�P�w{p��w>{s{�����#����_{������������s��So�q�\󹫯��/Y��5w���[�~j�mQ{|����~��/���wƏiGU����Q��\1]���{�ʉb�if�V�J-"m�NLQ����N�����$���[Ln�M|���,^��j֤�oC�f	�㶩gy��\h�q��(�4 �%�[�N܃����#?�=���ȏ�HI�f_<l�V�s�K�dF�8�� �9����.��L��j���7鷝�س���6	�\�l�����R�E��e���(��IY�5��Xȭ�H���P���Z�w�k�޻}EsŽ�w�=����W���˝��w��_���w����o�f�8�~�n����qjcutzx���z���YW�u�3N�{���g�y�����~����vo��=��`���a��P� .	��������6ᬠ� -S�t�
+
ΐ��E�t��愫�&\n|(�y�Wz��&�	�S)��s쑊�&C!�4작���A@3��]��k�p.b���&RDș�,E;y�k����YD_�a��������[+��	�Bg�a:��o��X�|����Ú��,�T�ﶝ�{W#�Q����gvg=럍mV��b#C�#%Ĺ���-nV�H(\r@"6HH�K�,$�	�A � !���(��8��z�;?�U�{U�zjz{v����'��������W��{Մ�q��ѣ���EO��VU�*ݒ\<�[Q@X\۵+���0CceB�W�3$I��Fl�ɭ���R��^>*gO$���hddf�HrE�M.~�o��^�i[�Z�<���e�I����C�4;�,5�'���Q���PF���=�1.h�%�F������zh����XK"&t�@"/���m�_А��2�]Q}�MQGD�D���K/��E�W�ԡI���|$ȓ���(�>}:'�li	+l����Z#	�ॲ������Y,��PG�:]J��K�U�����}��j�zA�H��G����9�`�$�'P">t�P�lI��,(ݢ�IS�lH��Z�u%�S�oBu������ f=[ȹ�S�/|���$���ρ4�'��0f`�`R�TSHÅL�D�Jq����+6� A��D5����cB`�I�U+sY��(�y
ucB��\g�h$u� �WR��P?*�a�@�u��4;��9�� C$	3C��^;���`�Z%��P��,������/�B�Ӊ�}�a�t�~�!_��gb�'$�F3>DqUg��_��A�����&w|����'o"�$9�h�$LsT_Ɂ%D$�^z]�*��"��(Ġ��_v�����Q�#�:}#$e,[tLB{}�b��%�*IȾ�M������E�/LH��.\ )�����bJ2�?n&ѿ�8y<N�Z�
FNC[5-������a(u��E���8��x�ep�U_D�i(�Lڭh7Ƞ�3&l��ք�d�����R�cf�"�����+�2�5;���J���\]F�垅��sd��}�Z�_�����>Ń%�$�~�,|H���r#h#m�&�N��0�=�a��!,w;$5�ݭ6�+vOKܓZ�:$�:zx=P�g%�Ǘ�}&�!����Ɨ:'�Dj؝4���Ȉ$A$Q�u�e��qHڤ�݈o�l���y�}Q�j���^)�|1P�on���߈�I�e�쓳��`t����Ե���$,���|���b���Z��w[O@��Z�yh�PYG�*k5qKP՜%7�&�/�<=l$L f�����%�Ђ���V��q�q�Pd��R�}x��5/H�x��$2�8k��*'����q�U�4v��đ�L7�V$0r��-$�����m�{�( �M5�����L
 M��TK����#�@�
LIe&h�բ(1^�ܶ����F`5;ٮw���}�Ң]�o��ە�k�B���ۤmc�7�� A��oޯG�_~~�?��'�~�����I��\��]�>Eg�S����Aq�A6��<B�R�����?�䓿y��W�R�UIU���O>��w~�R9�Jh4��.JH�>[�\A2t��Z����1�u�"�J�
͜K4��ƨ{�&p��S��њ{i�Φ�i�X��y��u�S6��T��>�|n���k��Xa������_-5��
�@�;���{(�=��r�F+�(6�.L��t|��͕�F�ïK(�I̋1���l��� ᓄOt�ٞn&zIz��z�[��F���|�z��I�4"�dgMs���o=����:���b<~c���v�>�0/���]��X�F��z��'2�2�vY�ב�2�% �,y��ƥ��:�.��y��2��WweŘ����M�Zv~�4e�KR�pz�!cf�f#0���s$L�������Ҷ���TM�r��)aI9S���U��(�߉9�7�@��E+�L���O�E��v��(kk������ҍ^D�Ϟ��Mb��r��e:ύ�|W�2K�A���H��<�*�&���bؿ
D�H��x�g���$���^�9�ƛ���H;m�MYzTe|�F(����d̝����a�bFf���ˉ¦҉��L��W"����N�)Cʖ�P�v)뤬���|�����+��|��׼������n�%�N���&Ν�;/B��N�|?љ�T��0c�����D����̩+� ����H��fLnI��&�Z�� (кo2� a����:�A������,�{���ܢ�����?>��S����떂}�������?|��Q�[z>N���1�b{�*5�!s2��*"R)j�'��b�~��v�Lc]���c���-�9q��'evQ;�w�~��V�LsI��/�'�hێ:��V �$cn:͊v_IG�<���V��� ww��(k$�A����3�aK������0Q�D7C=�τw���|��=�Û	mgV�/H)�LLL�=r��/���9v��ۈ�Bv�ң��S"b��hvi~�j�>[��x��1Wh"2C^��mA��r�1j�ʎs;�k�QG�H�K���F#�褶p�ɮ8�J^H֙�S�Ga��J������LKnE�|�2f�%�F$(�k;�e�ۦ��u��J��󗤺��-��k��i�Ӽ��n,ȵ�����p��E(�k�����b���;�Y�!`#��>�j v��|8ۯ��Q&�o$��h�Qy�x+"7ȹ���Q�V�-�7���ܾ}��<v��^x�O6���[�OO+��'��F-�}�+s_�K��h7�<"d<�2U�*�@sM7\(�y%�:�� �I��u��I�ܑq���KA�+!gn�������a�0k܆�]L�2W�Z/��Z9�K[F�Y� ʮGm��	[� 8|]e��i:�U}�ݟ��M���r���3�C|��Q�r�5�g:�	�`^DѲ��(��qeTF��
ɭ����$���x��M�<@�ve���o�t	ig�.�Yv����B�le/珅�k{֑Վ�g^q�U,4���E�:W\_��5�z��}tٟ�A��Y�.��o��Q���j�\~�#���FGG[��M��?}�����O�����_߿�={���=�3]x�[7��g�V}��lt����X��iV������{Դԉ�d�ⱝòt����p�t�)T1PqUe��E.�a�P�]>�9]h��k�/����IRvS�	\�)��C	Fl4��}���FSm��n�.5,����r v��͐�� �1-@�7����/
	�Ur%��@q���r!��mvg�င���+���(p\d�G"�*V<�Q4�rҍ8m����92r�Y9��t<����y�N�8�nvS;�l]�#|����,;?x�F�V�یu�a�y���=����x	ҫ�j��c�=V�8r !G%�T$�2���E\D:DR�}^�х��l��,�����7H�������;S>*��r�A�%��|W�D����D��D�8�@����^x�"�v�DĘW�	Mb@�}�����d���Í�{n�̙3l��>�R���f�:���7>UK㥆N�D'�v3*V:IAք&E��ɉ�<�D�I�0�x9j�Q��	���$uǪ�y�J����ߝ9>=���٩)�N�T��s��_a��W���T~�����ۋ���v��N��u��g�u���Y�_��SǻuuvV�LN�=V�KH��5���|���LMIv�<:=][����L��Z;Sz)br9fzeX�>���
i�d/٘�Sc�gV�G��2�>g�k$�s�ߥ\Xے�8M!���Gؿh;� a?�}��ӄNT���+�J�b8�D������_����x��x��ָ�����C�ML�����Ǒ,�-c��Eh7@�}�СCOMM̓���AE��y7HV��z��M
RfN��Q�^�a���9�_fl�������M�k6��l�������~���͙����by�w�N�=i٨2]��S�ɖ��,�-���I��2�!&3���]#��X�ZjT�� ���Qm��e5��"������A�w�n���V�&z?������20��(����k�g��Z���R%�@����Oq�ʝ8��@r���
�U����0^,I_(��r6 �
��Iv�����;w�Lϟ?��8q������4<��U���v�h6Z���.^�����{wף�0ȵ�H�E%��@0�SβD#Y%ZF�8 	��L'@2F���r�w�Q���Z����DfQǑ�*"IϦ�OQT�<C:��O
�Y����R)k'i�J�T"ɡd�h4�������������{�l	oA=s����W���.�-����إ��y%޶��l~����6ν��<y�d>�1	�t�Az�F �-�	V?�kl�0ξue���NS���N׽�� �7`+ ���V��V�]�q������e�!k ����v��Į�I�ㅙ[���/�����!��������GD��F���w���p0�UL��:�;I���ή
׶/r�'��ga�dgaa�llafbbj�p8�R��hN��҄��


	*2.,B|J�?���m�X0g�?x����sJh PK   �|�X�B'�  �  /   images/39b1e261-4cc5-4406-9e56-f0681178eaba.png�e�PNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  'IDATx��]x����l׮$�[rǽ�^0%q0!&�}�!�|�vw��r�]
�$�~w�gCb.p@H�Ā!6���&.ro�eK�$���e�7��٢�-y������̿�{�������4��"$��踆!AQ1)��A�4(�a��@3��ҠK��aּ^t~�A�����&p���w�U����fSg�|E�XG���Fas"^D�󸺀q�u��^�_���04���/���n?���a�h��>�`9�f�psMPL&A��nƑf�az	BD1Q�E�W`
�PZo��U���	Q�`b��W�+ʉ(6�G*��q�h.8�:1�L�n�E���A��>��F_�7�GÌ��ab���g��A�5����V*�f�!��͇�](�:�2��us+_�d��"	����ӷ�p�n����y��`��0G�b|m�Nƿ��1�8�M�1�	��l���̝gwO:�l:?��U�R�<��<u��0��ysc� ,�63N-�"�U��%B��B���֯V_p-I���صa"�-i�$����@�։�V��:���iu�-fe�a"ؿ��::Wa�$��~�<�:�h凌��s��J M���Ŵ�����u�^#���Dփ�KTR=�Nxrpuy�B.� ��k�M��2r��pXPr���t��H��� ��|�l�$[�
�� -^>���K����͜BW�'B����$�f��=\�Zx#}�6^���c\��:��"�y-O�uey���dx�S��-���+�=�����e4���UQӆ�œ�[䢦���o"vuq2��	��Ĥ��im��PW���rj甋��S�;�x����¼��_�c�۳��i���`���@$�ۃ�;�q`�l��fb�HԪF>��/�M�	��S4O�.t'p�@�A�ӟ#�N�Zm�f$�aqZ�_��e3T?��A���1hx�8�py}ݗ҆�h�WY]��;'87B��b�M�j�̵�]��R'��&�KbnڱF�}D���٬:s��(NgB��s��|[��HUӌ
!g�=��Z%W
�sK�����2a���F����/ƙ�<��,/�a�؅��l� ʉ3_�UC���ZH+�?�%�9zL���="�A�4��b��?�BNi���6+��"w���:�Ľ99�L%s;`��.���d�˖�q����i3�s��e�X�!���Y̪�M�j�&�)�P���N%�\�&#G ��	6��D�ZZ���6��:�����ط��bֹ�@-/�e�\�w��:4-"l���R��ַx}������;Gd�,���b���C�_L�e5H��m}99D#�d�0A�PϏ6��m�ݸ�:���qW'�c���Ɩ^7��GX�{	�#�CC��q�2Labt��ό�h!��z(!D��烙D��&o3^�7s��	�"��/�+v������,K���ނ\�R���`ơ��%�a7K �i�۷-H��w�mtmˤB�|�I�ĸ_A$@&��g��c�?����v���	|��j���A9C#f�^��h<v�t!���s�iD�"�׈��۰x�'����bTA3@�p�5�{I@�D�@&�3� �$�jH^��W���Ye(n��X�C�v���i�K�ey�F=��o����Oߴ��J �����`��e���I�v�������8@^|�����3JN��&��q9WE>���H!�)5�lbIa��"_�"}�Q���Z>�A
At�HA���gt��`���<i\]Vh��C&ܞ'�a����Kqk�Ȅ`���;HD#�3)�b��"7�`N���|'YW��pЪ�����1�]Q�fj�Q�}:^��^���H�0W0H���g�������|��I��6�C>nlϖkAG/rz�+u�&�X�϶�3�1���ys�����3�f��rēsœO7_�D+9���b����x^�[7%�������~���5t8n31X���_�I.20.}��s�I^�����BVq�*�M���q?�n�1sb�T�)G-�>�'���=>ɩ�ӷH!���,�v��O�:IJ��N�h�ɥ�lTDº�g�Ȋ
�7�0QM��C�5d�dD�:�x�H6�����8F�9���.8H��Ӹi�F:�����n��H��=<����C-.F��1�<^46b!�j�ܪ0UT x�tj<&V�Z3R��	��a���Ĉ����ܒiH�豿� ~�%�9GZ��ӧ�ۺŏn@��?E���>�����D���3�+W�}�dj΃���jaA�B?.��DF�輦%��!���$��,F,!��;�Eν���/Kl+�Ga��G�����_AM$���C��}�C��
$F!�H +h�ʍ�Ȓ�<9,���r����-�(����/�P���6<��﫯I�#1H:�s
͋���¶Xѻ�1�m||С8��\bԗ���ʥ(�4���'V�O�X3'n����r�f/�r�?R�r�� ��`j��}���Z<E"�V�9�q�nr9s�� �0O)��U��5��B����P�B9:�k����
~�-�+�PN`�:�c\F�Yݺ�5�-[r�(��ۄ|���.�Ժ�
�b�w�d�����M�A#������\�p���+�"U�N���e�J�_]�r����P�2����"�_�+vc��u�_��"�=��B9n!����B�EER�00�Ób�5�?/=[m\+2�����r<����K���d��b<L�IG�)��	bj���.�2��$�d%YA�D����$!�J3o����ֳg�UWcT������W��ىe��4�}5~OY](�����EO~^��Ѝ����T{��^)��,�\�vK�Qoi)����Ţ�;(�����-�3��>3��~� !~�VUm���Ί<珦��M��up�"�^K4��Ţ{��F���+C��Y[(��Lhh�;w'�-����KzЇ�5��+�~"��K\;du��xIK�|��!�N�!�z�LzT46a~{'�1+I�q1؜��P.&���^!�'A�Uum�ͯ �s���p/�gY&L=[���n0�4&
���/� ִy����
�ҚT߀`t^a⚢����1Q(ǫ�uHyӅ��V�<���'��d����-�k�"�a0���)��-r�z��r����āe�ġ�8�����2'���X���YFE�ܒ�v��/;n���r�(C����"+d�%�N|��<F�W�z{`=z�r��=	_�v���U5�}�*ḕ&��V擙Y4�e�*���1���0��5j�r�����c�эf����Ũ�5C���r��ʾ���h.��υk���^JsZr�� :q
���fK�}-�B9>ߕ��#�'����U�@ٻ� O��h�P�`��bu��(�*fs��w4
�r|�������<����]^^̠�Z��~�}�X����-2�9eq���3-�%�Ȓ�G�����47##@D�GRT�:����hh��Sa�X�Ph���hʱ8?���ܘ\4�������	�y����E�"K�-����~�4���`I��hʱh�R[���iKR�]��ޞ�y^���D�@��$��P0�rZ Ƚď�v�߀��M �5*2�����F!�_�(C�F�S(�ET� �+��`:?��ʱh89w��R�!de���� ���Kї��T׀;6oI�؇S(���h��P��
���XI�ڳ7%bko���C��[B2��Y����k�S(��B9jO���,��D���(�3(�� �D��	�E�����r,�N̛��7�N���֜���d�$�޾n����!�h����^K�t�rYS�>7���6�����ږ��!����^�5� � 0A�zzn3
�d�M�1[Y��py^���'��K:7؜��P�������ТkEL�'ARUW��W�	�yX�ڬ�����6��殁#�c�P���F+KU�����q�(��^��x�7����92�xb�$�y*����{`]�QY÷���de���CJ�Q3}j���~�iR�Je%2̱�����S&��!���������B9&HGQ!��%)fom�( �ⲭ��M����Vm��M��r\<W�=�)%��;��3�C��C�CV��-��/�S�y���SB'�m$��.o�!>/�K��R�.+Kȇ8�L�����P���RV�}+��Y��	�y��>2�ñ�j���d��� ė'�6�8��;�)ܥ��g��C���U��)�����`H��2�OԲ��C�v����i��Y_('ä	�v�{
�����=�L�T.._�1Bs���Y���V�d;ʱ(����S�S[[����XJ�S�<��}�1��Od\W7WI8�9�^��$��������|�A�!پ�[V\!����)VVM�9�Ͽ��r@l,s����X(�U�k�l�(Y���$u�^��М�Q���!���A�6�E��m#��o��p�[���)�1�N
:�~��!k�r�d5{�F`�ZA��%AdY���V�Ξ�7�Q�����p=B����"k)����c���H~l(r�M�˾�sI���9t�OL���C�$����u�,h���F�g?���J٥.D�������Q�X �
��^�m�`֬�Y�(ٱ��^�Kc��(G����yFY�+V[�wX�Ǝr��z����!�w�#�ͻ���"/6-��=:N��c����"	j(��q���c1�"������Q�7-.+C�W�����2ܿ��(piG
\��uS�8C�W��~|�����[[J^42�c�<��^�n}_y#s#��V�ri�47M���keێpH;�g:�򊥐,SI��im���y�`iV�Eo8��߃���:�c�ґ���s��~�Z�gLG��9���ۻ�%�0�����m\�y@����������'����G����+W�~�������7��������������!fn��Zg'�7ވ��&�S������G��1x�.!H{܏?�V�fw�?V\,����Ъ6U��/<t�Ç���G�/�9��[oE��~q���u��hD@)|&#>�܌��۵�����@���)v���X-����wz�}�#G�w�+��<~����F�	�<�[�����ۛ�@��P�cAQN�[��~�S�&OB�O \[+i�����E��r�.�Ղq�����{o���2Xfώ���o Uy���B!n�8�o��p}�s�5�͛�}�Zx�x����G���-[�7Nt{d�g�B`�~�3�q�čv!~��W�V(�:�n,羿C�d���MPǍC޷�%�����~/HTb;T�x��v�������q�i�w�{������y<��y�o��q?��8{�b�Om�}���> �*p� �| ��}J6��E�s�TY���>�ܯU8'r��Y��{m+���p=������Z�-ͳ�P��B�׿&���{�%8rD_�p�i|y�����X^U�s��O���h�myU�b�	76¿�M8>�AX��!d�_F̽p=�w}�� �׭��X���ce�͐��'{�������������"NV	�dG�s�x������a]��y�RbS��:]p������y�އ"���ĵ@���c�+��t���	(��B��Wp���~��o�c� d�0�������R�V#��o�q��\�mxT�y�̕�3e����֭�!�i�S(�'�J��p2�	��;�� �ѡ��<i�@!Nb���X�z�-m��bFX�F��VYO|=sQ�\�O�z#~�L]�OmB'N�qZ�=��fv�E�Ѐ@绿��(t&����'�z:D0a�s��q�b�c���G��8�7ap>c���Q(7��z�cQȌ|��9�_�2�h�|^�=�w1F V�"n�w��'�._&�=H�:&����nn�׉����L_#VϮB9���mA왳��ʒ-�0y�lR�eG��c~C4��;�'�E+9���N)�|�5TV�ed]x��	�y[�}��U�3Q9��c1�M�㩏&��m?Ώ~���71s/5x�E�r]��\����o~K�O��[���b��w��ŋ�~�IyÎi�4�"y��g�>�x_~��b�(���$�y�\r ���p~���+���[��bE��>8���rJ��+�Yloۻiy�΁o��Z�����e#��W��,#�������""Zu_��#�u<N�}�7����Ǟ�e�|��Do�--�9����f�ȲB9�a�b|����y���}�\z���MV�aG-��k��m]�BՉ�b�1�����,]J"�E��!3y���o��~+��+`�:EVT�5#!���P.B7��$�����8!�e��W�%����F��3"d�1���`!1��^��b�}�D�:�+�ǏK���z�����쑱-��"f6y��]����볳Pn87�ʟ��g�+g�/�h剏�r��=n9��~:n�*1����jB�w����q}!1�^ج~0��rlR�Y	]�-�vf_,�nȏ(��P.V�H���mX��
f�?mH`(P��X���2"�M��g���[���mل�������a҉F�i���:�C�/RƱB�~\��qv��B��hN���-B1[`*+�/'���:���]�j�V�(J��7V�(�D�{�f����*v5����:ѽ�(��/0��/���1!2qb����\3ǁ
6�׭�$(f�ӱR�
�=�'��W��W��\A���+�������    IEND�B`�PK   �|�XhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   �|�X�t� -* /   images/7a134b18-aa7a-4645-8200-8100c2fd668b.pngĻw8���C��|[��T[�����؛��j�ث�k�MD�ش�%%B�Mc�=�'i�>�}��>7m$g��{�ޯ�����
�A�@NBBrCA��&		��;w�
��/��\��.���/��柁��9�뻐���N���j��|H�Ճi9X��_;CI������m\�^;B��-S�$HH�(�|�푺2�jM�;_N5���2Ŏ�UA��[<\�������ñt�oV4"b4�s�b����=��爇�!?P��\e�"��'�6��\�x�]=
��ģ�
I;j0�7ig��uuO�A.�-z
�6��(6�&��r�9��L:�����3+��I<.H����i�o�R��\����%���5�#�����s�{��ØX��B#�g��Q��������H���
��;.�$�_G��C8׎��(��7�c"�����i��q�(\��HvZ��Yœ�Q{�*����:�7�V��qlO���~/ڲ�������@���F�?��N����#Q��K�G����-(OZ�N
�.����|�r%�L�>Q�'���%/Ys�;Ja�K�&��<Xԋ���I�r�q} �:��	��#&�͘p�i�|Uع3���궠L����8�����ˌ����~�K{\�!8��'���1���F?���%��t��3(G�!͠Y��-���d�&k��,O"X\G�g���j�^�9Q�)6$[�{fQ0NV����N����n�!�?�Hv�u�@*�т��@��Q?Lr���L\ڐ����p��%�� wm��,��X#��R�N�ߛ�V ��nT.�-j[ȉ�g~*�_���i��i�)g
�"X���5�s_B偡�7-�c��:2�9G����ގ7e�Y��=�s�{��a6�%r�2��@4�-%���`�ᗰ�k�J�5-ۜ�׈^�a�"B˰d��wZ�a���ośA�/�T<{��ʤ�3\��sc��y%��_�ǖ�Ol�݀�Y}�W�Vщ��n*�Oa�!��uKд����B֣BpԸy�$q*�.8Z�?�S3�*b��o%P�
��}��>�,
|�Y�z��ь��s2�6�;؉W��Ndɰ�) ˜^�J��P�p�AN� ���]0|��N����L��[�i�i��N9vU<�_�<��������IB�U��F������li|���oi�K��)j*���;�ZU6��V���e�`����:��������B��«��$*
�}��R�]��5:1�K��L�r斿SJ�8�r8m�]d�S�����KQ[���#H����p��2Q�}�!���f�Z�Hsnp��c{_v8�!�.��?���A��L(�G~��/�����#��s�c(�*m����&�H�ue��D'V�qz��|<s[����_{1�@�z:;���p_��@���IŘA�+Ӓx�}���r�7�!�o�a�EF�UG���-�j%�5�2~J��uT����_;�����:�uɬ�Z�^�'n��Ӭɚ��Ǡ�<�f4,*s*s?J��n��-��-�݋��[`�D!#�m����2�~��AV�|Ѵ�|�W���"�+��S�xyh�]��[	�/��T��.(���J�����=T���|�ފ���('	�%�nɇ5w��s������r���*̱|iso<��C3P��FM����n��(g���h���K'�ҋu"�t��`���O�p��ꓬ���JK���e{%�`��Tm	��� 0� ������s��?X,`���p��9���-�=��ݹn��r�a��{���NpK�ų��v;2,�p>��b�j*L�4�m7�{A�/�2�Ih<:��O�WF�i���A6Eմ���؀3hO�m�`g�8<�L�$�mF����kv�n�'̴�]5⧙oL\ڻ��[;�û�F�����K	�Z�!�Xɠ�꧀�ӟx��	>�2�Y�����
��|4��q4��9 	N7OpɶA&��-��^G�n��;8'����8��E�1��&����S�3���d}"B_�r� d��T�}9ӗ�z���꧞�}����Y����.%�f�|�s<�K��Lh�Lh7�C����[pڽ�6��G�f@�R�x}�ш5��NS��x�=�ݺ�aӠ��x��R���o���p&�״G�dJ���η<Fi]`Z��|0ߜ��)u@	��<�Y�������D���!��A0�n^[�� �\���ǐ嬺z��ຎ�.�Ro,�Qp�Mv�m��Uk��e�t����V��4c
�3f�xI#���o��F`4D#���Z�jO��Q�dDi?��ݙ�F�)q�T���Qq,[�]w�b��w2�"������3�^E]�%� �Yn�C_in�/伖��u]>T���e�9�t���vV6�ˡ���@sR�nK�:9�g���Q�r��V�	� ��M���5�
�^����O^D[FPm[Q��Nm�Ώ�"C����!�^KŴ��O��"ԁU�Q�x3t�m�������w�޷�ޱ���ɍڨ�I$-��I�&G�M\��2m�����v�ґ�6XX6x��z �H��q��;K;��P
�ZQ��w�c�-j2]�i����ChY�YΑ~#٤\�ٸ/��1�y�Ժ߰�߰�҆���y�~{`i���*�ݭ��^
���n�[�y�ԡ��!`� Ff��_\Dn�-�n���h�J����{��z)���<�ZtV�t��O�v��Y�W�!��*#��2��+���������ѻR6o�j�t�b�����I1�ܜ�ڨ�.Ю4��	Z�y�7T3K�l��I�����$7��Z�b���anS�Wl%�t)hJ�R�ŏ��=�AQ}��+�ʏ���x<�Cl�W�t!�z-�+�r/5!a���6�?�851�B?ἧ\6 E�,#�[���/0ʈ]��y%)�̖�:j����0�q�m���q�����w��~��p�(-�'�$Z0?��ͬR~�[4)���"0��	<16A���b*�j�����D��E����MG�BǷݑ�1��e%J��6��;�������ߠ��j/1BS�c,���n��"��25��c�YP��4���;��n���>d_�h��?وWu:�Յ8Y�h^-����Z�r����t�����?`���1��:�e��q�̇)��]�����ܧ��
�	;NCq��I��R��AY՞˿k��q%����axُ-�����d�4�0���^A�:���sgÉu��(f̧9w{��t]��]?+��2�#�ٕٓ�Z���C���ς��x�&FhLu�������4�w��^J���款s���v��C~i�Í��a�&$�a2&2tq� >]�,���󊾽I�)[��ɞ�lO�;����>�uI)�'$s�x���?/O>�>ݧjv ���7l-��M>JA�1���̚��:�|$�޽��an\sn',�ܼ�@���
�{��Ȉ�-N�{���ld ��c	R�M�V9.~��!��U[����&d,�_'FV���F<2�Wk8��V3������p��u8_b��n��;:O,"R�������:`��A�抲�NasJ������ʳ?q�&��L���N�Cl��шԺW�eݠ?��M���v�}o�V���gu;��.��;;��#����\78���+�J&q�\�_�\�H�t�,V�����f"��W(-���^
�D�z��@���37cB��)��?3*f�W���-�vո�4�v��-T|ڝ�����fgDڋR��}��'񹷷�%�S�`�M;{��'~Ţ-�ä���:Jx� �M����DFLl@r��L�=�u��)����VxE��f���ܘ����}>�CkI�7U��wR���ΩY*�B�������y���]ε'�F�u�Y�2���}WmDw�mG�갰x���=�w
V���aovqW���U����j{�ݤ��f���Tk^@��j�s?��Y��hւ�|�xL�1�$���B��P�����Iq[���Y�7��u���Ύ� ��X���:[������M��l]�[��6�Z�7�7-��I΢�f�ی�BM�j�y-C	��;����e�*�F�܋[g+�$�_Z6���2�s�E���^�b�N߶��f���3��?]1�œ�q�h�W��cF܀U>���}�X�k/���σ�:j�Ƈ6��HTS��AzO��Kj9����� �/���y���/�`�{���vbl��c�`�0�h}]81m�_��y�>E�Ѱ�3���޿a9�؜t�mr��/Y�n1��T��t{_~̋۾��^�� �(�]eϩ-Ƿ�1@*������9�D�⾏��@Q����~���6���R���6�:�:g6�[�Jcc�=L��O�_ҭ[R��cO)RA?V�S���[ZY��{j��B-�7Z��o�l� �`W�;��g��.�-k��|���M5�ۛ���2&�AJ�i�%M�}�Y���Ӯ�P�������]�\�`vL'õ��Lp���4�@PPBx��	��U<2[�J�TAo�t�Vy`� &~��iy���GbL�Z���&�@E��)���s��D��s����y]*����D�(��.����5T>09n"촑�W;�[o!��k-�y��U9h����Ц�Rt)BimE�2� �|h9�η���W��49��SXlQ�W�9��~�-�\_�����s����&�#�����0�z�T(�ո�+a9�hJ��F�p�\��;�R~�]�D���t6�ڿ�<��|b^��aO�Z�w��5Dz�
��k�t�1�|X�$Xk��~�Ө{�����Z�@Z�'�f��u	�p�6e)אYB�i�u7�6aS/���`��[(��=��fj�O�An��yr)�PM��r��|�������Zs��6���T7�D�5���Ǧ��z���f
mq?� [~�h���] �5TN���}���(M���|���؝�
~�{��ֻ�,�z��� v���V�]���O;]5��ԫq��~9^rJ-��;-kV0_����ޤ	�M���Y���G�a���)��{�z���WR� �1�ևk��?�]�3��s���Yk9oZ5U^�`�
�r����oh��#�]�e����mA�_3�� ȣ�B]8t%Z���
�*�#E� yH��}��Cu)i�4hp�s*罣I蒜��|:Y/��O�� $;3�݌Y -�w�~�D��@�u@S]%EY�2/���Wӵ�6�8Ê����m7mqAAACa	�
���$���S���%^��;٥�@˨��Ƒ���.)4{W10��.��V�O{�OKe��Ʈ8��&#���a�����ӊ3JѺK4�NO' ����#���)���/:�z�h ����ig�y^J�=���lE�,�b�I~�E�,hZ���-���m�d�7���Cl��d�0�А����Џ�y-�.�a-��B�7�7%��4-��N����$6�a���� �X�1$z��8��J/.�G�$}���x�ֶ��a�K���Ij���:	�/*���A/8��i�%�N�0b��{���Q�I�U'�z��|����D���I�_G6����r��(������dm��y??1��+>�f�1��`c��}��n��Y�Yzh���4���Ӣ���NI�Q�����ρ �Ǿ�)�E�w'�j�_��:�|US��F@=+�x�����;��<VɌ��uAS��ߗ艺�d�5�l����}�t��TCY�^F��*�;�so���[�H	:�Lˊ5���
�P�䦧�W�=Q����\$g�5=���W�_>�]�O
���&wW��f����B+[r����Q�9DTJ�-���.m8
୊o�6�U,7n��(�s�^���Vf4�ϰ���9�����KV���t�L�AD��~��8�"�l��8�Э���Xn9�2�0Lp�8�rn>��1��S��'�ڧ\R�@��}>�t�� �b�� �����,PS��`娳q<xA=�vm�E�}r��f��`���Ҿ+u͋�znd+ه՚Kؗڶ8=�Mz�P�=�{FX���i�Q�QPL��W�6e`�A��Ў�Os�W~�!+��-"CE�;P�]b�.�Ͳ�ż3��U��e\C�N6�Z.0Y���t��$����~I�r�p�L� �|�N�Z���'b"�A��yRZN9~G��t0:w�qFb�Hk��{8!�]���9.+ЇG#v=��H��ҥ��9B����k�j�O�u��O;��#T,9d�L�S˙"l�������0�0�B|6�L�P�E�����h֢y�%	��=�̙э��������0ɞ�S���.��$��R����s���c�I�o��5��L�߈IC,ߚA�@(���J�5����|k���6���yl�S4	Z�؅�?U;��K�g�P?�D�4�Ǚ������p�+����+ Z�~��!��w�@�UoĆMVw ����ol��� h@�+@���>\e��S��|��0���gq�&LO�6��Be���?\���kr�8��1�1�h�p�w��< jhfXӽ���7���Є8����\��c�>ғ*�^�Ax�<V�4{ c��T �%����X�ل$��+"���wjq
b�/��?t	� ��֤����o`M��Nx�(��l�e��?�jl ^畓�ǀo�lƮ�\��mYj8�G�o	Nh�5�3�,��(}d�f����/S�]���Z[B `���/]\_̝���X�krК�����~��M����Y��� ���������낱�'��a�Pqm�MbR��S��hm�e��L���]b?�7��;�F��+Q�qG��RG-#֨��b�*����� v��Υ�3m������Kew�{^;��U'���E�M� ACC�fPJ; ������ V���%@���P��'�C�yx�dXL�� X7��E.������o��ǚ�ޑ���{י�%x3�:���;�#�ڨ�D�زn74�Z�ߙ�j�f��~�����E�2�0=8
�5�	�9NȉP�
H>����	|�ux6�R���&}QﯫB$bV��f�l�F�.p3��ڷ��<R6\����k����"M|�dL�B��m��}z��z��	i�ޣ�9�<��)�Zd7(�4.� j�[�Y�4���-x��)�ȏoT�cv$^3*�!h5G;TO��1oP����="l��M:*�%/�Wz͟�/��ۢh�ȬS��Ǵ"�Nv%� -��4,@�)��X��j��ۤ����;6%~8ߡd�ʝ1��^ݰ��1���+|�5̹��Y#����E�=��Hf��cj�y���D��Rַc2���Ø�hJ��$��|�o����e���^
�<�δ�aa�e>��Y��X���p|���͇�eۦ �+�Լ8
 �ᾌ���A�3|�]��K��~�طJ`�?�z&�
����|�]
�񜛗���Ų��d���
X �4d���� O�����0��jw�5��t|�u`r.�S���2��Ѐξ ,��~�\:3]Ii�>v]-D'��6��?��*(����<����{1,y~��� ��=�m� �N��x(Wg�Cy%�x��+�gR�℮�D���O���g�,�(E���瞧��g��ɂ]��oA�S���	��P��O�G�Fw�VrǞ��$L���n�QR�Y5� �H�x	K]����t��\��Ḫ�d�wr6i�"���E��wQ��:4�(�����aZ���u���ۍj��O����� }���uwU�-e��,9+].��W Փ�?�n� u���l�;ҺQ�mU��:]�ɒ����|��<d�q�����M�?�ҫy5�q�����m�*��γ��'o�c¦tvW�r$� o�L�����5�t�צ7�-&�����&����ָȣ��L�J���P�i��q��u����i�s�u��*�!�X���x����/���-^�(ܯ�DLyj���>rfL���k`�����J{K�� �P��K����/^$�A㡽-�rhnNtF���w�NRo4����t���x����Ŵ]��E�53��?R���m������q&_*c�z<O�NǤ�@����������f]��,"58�/m�X8�	Q�<㟼/��\�]s�^��D0�-�^�Vܣ��r(B`	O{��j��5��>�H d>��OafW�z��;�1�^��7���
�\7�6�5T�7��K�:�W'�}����]#�ȉӟ�����NҖ�$�qz�����֛@�����Dj�S��D��t�v�I���#���!ӣ����k���f�wRE�{���$�h�-�p�ȡ��[͇���'�v�=����|II��FͿ��>�W�~�oR���W�s����Ze�*��+�5������wt^,��Yx�qOD�^��4�v�񣍋��2�?p�p(Q���U�ѱ��8��컜�!�6/_��ٚ���^��;i�<�_���j�J��-f�e�Ji�����p�';�_,��P��K�R94�21��NN�Jz��j��5���qLKf��LHf�Kځ��."�(d�����6�&��5�h2��Dj��6r���a��}�FU9p�;�鳋<�^��w׊MA_��0�CMr�NM����Cqb+�r���,��Euc��ԙ�N��ube]�_������r��v�<?J�*C�v��RQk���a���� �ٜ��	Yj�'p�Q)�"5���DgȻFw���DO���!�=֓�S���.���4v"N�����K�� V၄��~����n��`���}�֏��!��._M��E�����:{��,���W���X�8-d�9z��,��7Q�gb	R�O�G R�G��3��%�I�;��}��!���I׶�7Uq��F�ߴ�-k����+�wϚ�rt"W��,K���xT*+�Pړ.��'w��&N�~f��F�A�u�� �%.�D���%J��"�Q�\_����X����CS�����QG�G	g�1�C]�%�\��,Y)s�>�t:���䮓=׶�ck�'�wk��DƜ��I��f�^�j���%����΅%�����Q�u�ŬFW�o����$�1��$J�1���>�����cݚ��[�!�J�|���d8�ɵ��AyMQaA(N�a�-����� �Kea�*fz��҅C�̻��i��փh7LE��a�:c���?W�8�����fJцy���l��Y��B�kT�p]G���
�����ݖ��>�m�ɭAw����[\���.CȢ�d%��[��vp����v�i�-ao.Ɵ��M:V���*�<L�0b�{�
o��zH2zܿY�����g!�~"�8OEB`A3.�.�2��W}ٲ���?�˰����8����(���дRO
��~Q] !��V� u/#�
��ӽ�&||��P�{����aW���Ct��wTsU1]Ҽ�i�GV�Cù������r3g�SDÑ
�x�f�Q�#��L~�d"�Lp�F�tv���8����c�J^:�)/�N[���a�À���2v���IS��D+<g��!v8�Hl��NA\Ue<}P�>hIƔ��6�V�#��j�����z�o<�j���n�XL�[Y���K���������_�:~�����D%P�s��2�~6L<w`�~4^��jMi׌�v�!)S&���0+Щ3�1�O�:*!b�H���8 _ ړĺ��<�����H.�a"�o��nP���]��6Ư��=+EtE���Ҙt܌$��~�=������G����ֽ�`�����0�YCO�8v�ъ1]:*��H	�WQ�&��w��47i��!�O�_�2�4V6������� bH#U_`U�Ǔ���[��J��<'»�CPLƪ���{�s���P�9�b%�7��*�]�|�=we.d��o�C�NS�=�UȜއ@����`3e/�}n]��C6�E��n�	�@���hw�Z�t9��E�p�V�ub���6.wǩ�9�X�[ ��͚x���ՎI���'���������p��cp�+�6��w�>�HJ��	�d���x]�:zF�Zt�s^�_�ʍ�X�y��@ߥ�����^<Ц��@Nk�s�=�Nf%�7%Q_X��s�ևs	��x]���N��  lA-Rh[4��y��;fq�9�8�oZ-�!.���@����KAE6˙�	@��)*��d����ǃU)С�!T<�A8r+_��f9����T �g������_�Pw;� ��-��,��
���?ƭ��@�[�MH ��ꕺ�}E���,[�+4k���H���x���P�'�ܼ���{+Q�}��?���P`���d��� F6�/�2L�v
�'�r�SZ����^�%�t����>P�VD�>�D��C�&}� �O�PZt��+�Z��qOCA!��knw�0�"R#��] �7�%G��<��
f���'��A���]Q?PN�G�;s�ܱ�4��$u�~�&��-0�F���-ɜ��9N�?O��Gd
	�܈��->�W���"��0?�P��6��;B�涞�tv�K���$��k7���1A+�g�1���O�2�t%}2q[��;�#m�A8���`�]�ڥƴ�dԵ
fּD��;0�-bJ+�t�#��@���������B�]�h�+�Zk���Lv]2a�O?�c�M�r��A�=v���ӗ��.�cIj��@�%�?�g-��cv�^;5o	�D�	e"��8,׵'iP��ɲ4��"������zg�)&��J����8�z�IaX�����������H�5���=5��KR!?���}��V��l�sմ��7�of�-6u�G�;}ײ�����u��S-�2�`B�n��9��Y^�����U3��֣B O�r���ȱ���5q=y�j��gĈ�ޏ�ͨ�����U��Z�4�`�Z���U�E���ʢo�Q����4@��g#�� Ձ�]�}�1�oՠZ�{��sy�<bf��We'�$��E8/I������̋�Q��g���s6����s�D�M���k�?B�f=��b�#��̻�֫���"���>\f�ej+��L����/��!�H�lQ��)e���|�[�����0,��~����!Y%��<*��!HB紏��N�ɼz9�4�c٤h F�ji|=JH�t����V�5n�k������^�<澥T �I�R����ޫl��}��Ng�v'��߼�'g�Ͳ~D�D��f���w�:K @��� [K�}<*{�yǟӣ?غn?���\��RG�����Bo�ߪ�b"�����1􇳱�r0 �1mn^��S�������Y0p᪳u��Sb	�学Nl��sO��"�GT٩�hm�gI�	��L�C��_Jk�ʚ'�#R9�� 3��NC��1
�B��>�5Q�_��EΦ���Ł��~��;��Wȧ��-r�,�r[��:����Kj©�ňׄm��)qǝ���Mq��_|%�	�t֙�
,i�a����PA�Z֫L��5UO�s�K�L��^����Xc-3��g����.y�S�s�T�É�B*=�J�ʣ��q�G�]n��Lt��Y4�b5Hb���q7zގDɍ,��h���*�q�i�SC�'��V�V9r�!L��F�V�U.iE���E�4���TD!�˖��({2z��*Ǐp2�K���(�L�˦'op�����M��&xU�\J��&G\zᳺJ��	����͗�H�*,�u`D9��T/��.��0G��8�,�<
/�7��m"�K��	!l����tܿA܋,���C��w����Zg��	�k r
RG�.�0A�Ѓub�ɩZ=ʻ/��)H�N�u�0
��t܌�㷛� ��btBLdW.�I�+��
����A����f�4	І���+�@Y23J����"�q���:�6kg۳��8�c�#,��Z;mZ�����@��!��O5މ�u��B��s�%�~#���붜=�Vŗ�N�\�u�A1�r��m�-[d5t�vV�t�����+��+�S��2B+�!+>IŶ�4Wys�<ڰ|ڐ|�u�xus���Ԣ$�!PN��Q�E	���/�]��ߘ6O�h�L��]TT~������(�(���$�8�*m�h��W�}t�
C254�O��~�l4=[��H��`�d*�\��e����ff;t�b����\wß�[�`�����徿4���}Xv�I�P��0��R�CK�O=$MZpBO	>SM�Ym��Z�;S�=QM�rgʺg�,� 3;I�U��/�һ�4Mϱ�Wio7��4��2�����E��Y.�H)����Q׎���bt�%~ar��+?�r��Epx��)+`��4��H�e��#�׺��S��( �HJe"%����.�ޱ|��L��e#J���:�ٱ:��8�Z�1�-zǮ��@�0]���������� �J�
�P5~na �d�p��l!e��J���-)���I�Y�����^n�tE�[A�b0��A*��ovPR	�g���ỻ"���jI~rw U��R�8��^��7�@�*��Y���z桹����D��%��3�V{k��j�6��)r���ݻy�f߾*�E����L��v�I�7ӍBJV��^�H�8�_��Q[<.��!�c�ɼ�DK+�p ��~��<�z��gز/d}�E�o���V9º$�}��?��L��U�_�U<����P7OM�g�ߗ�
|G5{����d~"^ Z/��i:��i\��am����Z���Ѹo}v<� $b�I��O�ǔ���%�É��|1���4�囇�ӵ����ϵ0�$6w��YB�_D3%$,��l�S9_n.{M<�0�O�^m�TYW�#�DZR��<��rt����J����	��F�]�τ'�p%�\q7��(�YkF���Ѕ�C���I�!"���o�{"'�W�ߞ8�;a�w���=~1�Ǐ���<=�h���3�a�?��<�඾��:F~I-�M
�!‿j��1��'�2Z'�ݵ��|�E�2q��W�8�3�9�����l�j�|ǪiͭOfR������$�Ul��8)a/s�s�p:~}.��}�I�KFs|��z��_ڒ���9���Фa��걓�T!)��P�n�:�����>I���D����q����VI�[�w�t9`z���o�WϤ��nH���A��H?"w�w���HTdN+�M������>7�9��X�g�/�h�TlQ_%���m)&V8�!8���!us���7%���AR&�E7?�0��b|t��m��8� �����|��u��HDX4���.�-Ty�Ғw6��R�_�T"�D��E�ʇ�¥H_���T�꿆��kس�OC������F�٦����I��p.~g7yЮ!5�c.�p�p��7_Gx�N��ơz�����$ޝ��j�;~pn�����;�v9یlk>=@+�F���=��wl퓙�;�Q����3 ����n�8l�]��g��{�-�RͰ������gP��ñ��Lsh����l%v�=_L�ŭ�Fݎ��0ccqod�0#�ߒ7��&m��)�-���]$.4�5m�G)
&�j�0��/&���y;;�~���t�hbr��&��A��;��c1a��h&�\[��;�������pؑ���4lRWtJ�}
��u?.N&-�?-�?F�~�5�m&O�?�4�"��*��8��i4��L�����4r��"쬚�o���(��ŀŠK��'�vJ@���=�s慔ۉ���uG[��ޔ�a��f�Gr/O�����~�T�"����p��4ڊ��>`Q���%C�m��Q�c��q$�?6�����|t�����<`k}��r!��/����x��"'�N�ٌ$�(�[?�P��Ki�ޙ��nMʺ�ٮ^9� 9�9�&yO>M0��M%�msQ�[T���A�������"a��b���+��ꌴ�b���o����h��S��omo����d���B$'Cv4 �o�zSw�7#�$Ql�/�������Jq���%EFv��^a��O9�Ҧ�K|J/A0��"���k�J�H��	%�.����0���I,�������������؝̦��SE/����t�	�h!���Q��e<*"+�׍�#6"��ř%���h��=�l^!�˪��$En9�n���yn��#ڴd�����Z���m�n�Ĭk*�u����s�7���«p֣�t�����5@�[��1�A�����&�Q��
��^��`v���U&�N����q�,���D�F�4�T�-t��r[��n�/
~W\����.� sB��&$���N�,�!F�y
[x�@��lQ ���㴫$��FiRd`�b��8R rt{ao�����E��iNs��)�(���z�n��K���̹�O�z�
�,���E،~��w�����b��)r�-jȷH�7 UUϼэ�Py�Hӂ�e:�����h�@�e��a�� �k򺗫�u���V���bF$Ϋj�?PMo�@�T6���|e4q�'sj��eɸ��7�JP�������E�5�Fϧ���a��h��π�t����3D��Q��4RW1�R5��q'"��gH@���n��(��+�mn^�F+�4��CQ׭��}��9&T���㿘J��4q�h4���G�@&Cty'�M��Vdz:��F�����G��4���Ne��$$�+���}�6��
��N�ǹ��TO=�q�(����_��F޺�p��Se1�W���l?և{y;(MX
瑩3׫^w���rY8�C6>.����s�u�X��7��/�$v���5��Yཞ�~�ޫKc۟�����
���LZ�
8�s6C$ �6�3�F�O]�w���7��2F��Dm�ט�4 4�����H�H}��R�p)j�R��wYU����vr�'���%�6��6��@E��"��®(+�~$�����F<F.�v?��[�7�ǇCa�4>�J���1BpZRr��~�H7ơ��9G�-�W�(�H�2����ʃ��-6,���]D?�@5�#���".��pT����4�:����K��OeQ����#څ���3��FhϪ~��ë���, ���������wqm�JqGB��n��k��܂�F�П� �[IkP�MK���xs�k&��ct�K��uR���pw����#�}1����T+�}�k�Ô1_�ې�.��U�wD[����<���L��F�	3�Wj�?��j9���w3�ܬ.�%&�9�wW]��$R4CP��W�`{C��:�R/�n�⯷Zy�g�t���E����R���y�Z؜�i�������k��?�{��0
h�����3��=y"�\,\����K?��?��Ύ���쎽��8,	A���=����F3��U�]/�Z��
�.�nu����R�遛E �Rν(�'v�Qi��k>���ao��j����\����3�|��}ѿ7ڍq2K�J���(g� �̓��~��tq�"��2f��騧����d�'a����y�$�I����r�ҁ��^�^#�է�y'&R�������|���H�o@�����|�oT�n�66y�7����ێ�����g�"��$B��d�7O��O��9���+��ӥ�9��4G�;+�	�"��(�����S2����xt]�
��
�2���1�~�ǀ�x�;�Q�k��O$*_*19�|H �_W8�W��XX؇���RTM3?���$i��T��п'�O�w�j�D��	{�_ݐ�9R܆*h�5�r��U�1s����ⷸ�y�g�����H:���,"��B�"i wz��(j�
���l��D���R�U�����y�0�z��������f��Z�۽F�nw���2�e�"Ee0�	h���F�_4�J���f�2�o����G��RI����sO��\&�N��]y"}��0��eW&x��R�I&�^7h�Я��Ci�&E\�����UMq�[ f�����I���2	��Vh����A��b8�Y5)>��P�4<X��Lj{Y��=��Z&���0z��A���"�/������z���eeC�T����i�B;R�����B�{rͿ�+�Pk8�X��+�n	U7�DQ�v�2��|�JaG�����T{Yb�{TM��U%��@����Zy�uz�l�M6l�Sq�d��d,�MS��?o��6rJX��#᪒�����׻�#��q�1[ڏ����+�����<�5n��4�'�ث5��������r\.�,��=Vy��J%�s/ԭ��Ť��@\��?��E���945ހ���)�J�E�e�Hb˶6�"�����q�@N#�!�W�����+O�%=<i4�|j�Oǎ�-��vC_��ە���4k��pɂU[�/b������^58����P~��eNQ7��ⴌ{��~�ϦEKL�{��D��nB���;�,E-�(�y���"O��yq�%p���#�n0�]��=[�Ӿ�󍴳����[�(Ƴ����g���!�Q��g�8,nZ�]�I��fXP����	1Z7�q�E��c�٩b#�`%�Y����Ô��M������z��C��*���K�i8�WŦ���LSCӡB�ȕ�/c�Jf+��Ͳ��L���3�:�������7�>dV��B'��)��FN���{�r���o6��%;b/~���8R�PQ"\P��t�y�ʫ��^ S)�n��o�����5����*ՙ��� ���͏u!���L�(���f"˷�ňA�t���3��2F�V
�݌l�.�>}�Pz�9w�έ�(���)�HD��i�Ԁ�7��Jm���.��s�H��Y���b�"4*d��]��bF��4��^�͡�����q�y���]��&](H�̉G)E59�n�/'�$���#G���dMo��zga�U�ɳ��.z��A~���F�-3�8�D�u�_2h�����'2TRD�mI�%��7 � ����-7t�{�Ӏ��,[�B�&��H��
���/�RӌsGD�|3A,�8t�u+9t��b_�tF�Je�n)U��F��&����Tu\�e�����+��UQ9r��V閆�<HwwH;tw�H% 5tw#H� Cw:�tq���u��|.]�%{?���{?���z�B���S�w���{�(['6pO�Ԝ(�{'���"T��{[ 	�o3�LE�;����������1��χ̘��Pv\�f��5�������>i�fb�@�z[�����҃i�M�c�*_�`v�=F�Oi-�����5+O$JO��kw�Κw�6��U���'�F��ݦ�����@�͵n� z!�9YQk+�MO(��t`��Y���b���
sɁ5��X��V��LS��N:�#(	l�\M��H��R��b
�26כ�	o�r��cK�=��֬m}0߸�(�yܒ���M����jR��_R�?��ޜHz8�<%��t�5��.0q����8wҵI��F��걠�Gi�B�S 1�6�uH�C_Y��aWϿ;:�� �Յo]�;�44��K�}�8
���b��R��[|El7�:�y!w�����6E�8������,��Hd��ۿ�+�{f�/^���+r�EFה����4�u���ΛqKk��%P��S�K��]]@9�]�.;0���N�e�I�PѺ�������4]>>sPĦ�H�j�,B���c_�z$�VJԢ��9V��au��4���u_ܱ��q����(�d���A�/\��m'�Ť�1jk��fz��������7rE8��t����V'<~Go�*_����@&�^�A����Q:�m��`�^�b��o�������:�X	��oR)0[(3�ױV�'�e{�G�����t�4z�(��������ę.�)("5����W� U�3��D�?�Y?��t�����;*;ߩ�C&7�c��8��Ċ �4����`�"��a
)B)}��y;Yx�]��>�/|�1�*�$�۷Hͪ�$ίj�m_�` ��.��7��嬯v���v`�\i��ƞ���:GQ/�t7Ek�" ��B�fB�9�����TҋP���P�9#������/���[~�B]� }S�Jc��(�����?�:�u"���6�sלe�=�htCk��a:j�n��1�
���Î^�^k��m ���z�=jZ�2�oD5�?��O�G���anS	*т��k�c;�*��>Z�ZС����r{\��[���Iz�	�Y�3nx�)U�I�g7wSa���F��E=T���m�,��}�r� �J����X�)0S��ޅ�EY0(����k_ic �@�� ���|?"=������4·xNڒoR�y�h��A���� ��Y�Uw�m(�F���	\��8���v��s�P�Z���W���GP�	�]�~�;��io?#�O����O�	�8@r���K\_�yk��z �Ԅ/�������_���W��A��M[�S�E{QE�˰ <��|=`w�3C aRVB��[�*���
3"νԨE�\uɂ�\h_n�w1%�Z��=ݴ�n��\�6MW�>0/���R�V�J�ä5,����]s�D�[����[��~�Ke�0�Lν�݋���}�P��a'�̕��.'�\�?����g�����Hʳ|��h�"� ��"'�{�Q!@��brg�Vc�m���G�M��Q��e���!�c�u��+�8H��●�9�d�X�>�O�= �e)]N긔���+�)��6�7,p���'�l�����C`E�x\L��8CG�/P@壅����2��TXL4�ٔ�<GFOZ�}�vY0�4f���̥�x���d���1�p�}u6�۾l�/ݛ���d�}�A�b�����֑����<c�!H-4���aɭ��?��H&G��aUgB��ń�S�?6ܥv/A^�Dck�Ԉ�Te,�  ��
�r	�,�K)X�!F��S��ц���{.K7mtl�?q���������������-F2k
�V$V�y���њ�N�u�[��W��A eӛ�c�V��i��U��|��J$ep{☧��S�(�y� �d��aA%'��)�PL�����97�=(4�n/�a�v D����0-����[�īWy+=��z��6l �D@��d�b��%FFF��:߁Y�<a �L�ĵ��X�@�
�?��
�%��<m�v�ēZ64O���$S�W���'&fk9�Ɨ���+���ӕ{]{۰GT��{/޵!�zȧ�ay�!f�[������r"�Z��u��Bm;۸�~h����^7�,����x�L��9��J'�a�l��){A��� �%�X�^��M���bQ�K�A����\���Z4���T
�e��I�����^��$�(�J�x�*�ǝ֩�t���OP��"�zvX>�"l���1��7o'U�
��5/���J�r��t٢~�9r����E���*�(��#�2����u�����ID���H<�XZ����m�n�u*�*]H��}��'G,�G�e�^-TQ�Ib��t�y�mr���t�o�b%���GKa.�П�$2�F���N"~d�}�<�8_Tڅ��i�ݺ;��R�l�r��������f���9b�b��h��oV0�Xw-nBԊC0^���h �� �UZ��In���m&&HWLמ^�����*�J�L���F�o���8����D��6ۀ��^�֒`9�=�4�N�����z~�ܽ�B��FX@�j� H��=V���s���+̱E�K�o�Ep�ؔ��VVyn��U��_G��i��G��z�H���F}��2�J��޽��A"���n�۔��ĊBEF&Ipt(�pLS�Jt�"`,�6� _�����W%��nL�U)����$��R&��5�_
8?�Bi��_��mll�'��d�$�]��E.`A�ھaZ�q~�g'$H�N� F.�HY�%�?| ��*��\��3� \S4�s�?ݤ}�iF/\0a����N�Z���C����E5�Y e�{�'��S�Yx�"kZ��- xf��o6��������!��J�)�'�D��vĜ�Ay���2��ZȘf�{,�{�S*���v��dU�v"t���u_��~��g�I�� �A�}�n�>^��R�K�]�^a"��p=�Y�Sֽ
3�O���I��ž$M�u̖�S�o7C�T���C��� G� �������_�=C�l'���ϭȆYq�Ri��Ӳ���˺���=�tӸI�E^.��e�,��DÅp~�9!�3˴k�}���(�@騄����_������L���+���"���5=4���rB�J�ߎ���E��p�E�V���a_w/�<D�կk ��t��hX�$� ���>|5S ���@�Ү��ϐo�� e��ӣ�n���()��W�rGa")����`j$���� [i����jV�#"!D=�,�CM��d��IfʁXO�}= ���?�T�q"v����ݛ�bv���D,A7鰌wg.;ix�h3��w��V��߫�A>��ę�-����PY�e?�x�ӆ���F:�����]����Mo�5Ad���M�~��n����� �/�I9@�r��I-^=���:
�������r����(@T��tL廤�T#$� trҷ�4����@��%R��.F��w����O߲��7n=+�~��C*n˹�v|���{����Iy��zvQ_TAal ڋ��˝�͞��!����mA�}���9g�/�C����++?�L��2~����B�z���䦥<oA�RFB��@J���2`h�:G�p����r�]���I<]����B*�w���o7uJq���m'��ᔭ�l����8���M��cƛ�J� 
a��׹\�7!GS-�����'�wn$0��֊,�`D;�Ы�| 7�gz��j��J��ʇ�Q���w�c�uJ��۴�r��{��o#�2��U�ZJ�D�:�*#�)q3�G[|�Q���C #�#0���^���J�,�}�ğܻ,��2�&Q�4J9��@��L*9`�*��oT���@��@�$!r()jQ�ֲ���ғ�j@��:4v��Ԇ�=���`!���e�-�����ѓ/}4��]��k"O2	od-��N��$3��7ق�!n |�Q}L��m@����`1;�g���4=WGM(�{mA�3���v2J���Rű��T���n�
6::�Ά}�H��i�lJ�b�֜������sϮ(J/"��n��g�h� �N �6��8�}k� �Ɣ�4�����!��%��t4�q�_�YM�s�;KͪҋW���֚<��@]�m2巇5nt�rY$���<fs�t{�V3�>ަ1�K3 
X&b��6�n���E���=H�c���$X�	�1c�ֺ�{�q1L3&j��  ���5�Զ�>l��#�&{kMwG�����F���{h@���Ba�mv�S-f�u�u�2�4�Tj�]b�m㙟�l�?���Q��&��P�y�L�U��D��	 5<u��e�tM�*�g�pVXV�����oTX�<��Sm����͗���г������|"uI���i�h(%G��)-���ڹW��n��-�-_��̡H��A
�N���sY�pfq�+�u�X�"F�/�g�hc�63m�>��9/U�v�(:�m���x��$��V�VoO�jD#��J�p� 6�K��O��� *0�2u�Uڪ�P��<��\���4ʎ&T��[���>g��v��5d�j���*
��=�t����a�,����cv�֤��I�p��F�	7��w�M��RT�9J��}�כ�j^�7�ڞn���	����3;Mm���H�\��NA5�"��xo��,�]���%��0-{ ����8��7�H����Ӝ�gg=''�-A
IuuH_iԷ�Hy�^�q��
�]ߪM����l)A�(#e���(��O�����z�׮�q�����'��OWg�c�1vd��<jԀ���-{�wMb@���@c�Z�\/\�9D�G[����빈L��|ls�� W�Ω�+���LX��۲��c�5���l�w���C�Xp�
�����E�h��3)�v
�V�|��;�.������d��"����pE�H�����g��CyZb��7��NJ��k���]� }ܛ��eJ���D�T�N�Y�a]}jWk�cn()��A4p��mk0<�òa����@��/v@;��f5���� )g���c��iD�\/~x{����#ڶ��[�ڲ�*E{$��M���0%��^�o����g�=��G�'d���hX���b��E��;g�s<FZW������*����L��[��&m�7p�Y�����l����ʑ���K7X�IqR�%����$涋�s��N����F�e����ߪ�L¦@�#c�WT^��9C��52�62:�͸�ט�%;3��D�����v����JO�2.�hz�j`�t�5�]�,$�9Z��`��H�̻�����2�
�T5���s#��?��w�&*]<��5��)*��T�\�\&��b "�h�L�IcN$Z-��g�Ha� y��|���|v����k��O�+��+$g�avh呏�U�g:�<(#=���q���Xl�xM�̮���������nIQ��l��V����T��@[�\�?(q�q%N�����F��妲r�!FF�F��R��2S��3�&��çD�eLa��G0�ߪ�	H&)�e�Ē����?�*�}=\P�vySL�t�mn�ɗQ����˞�I�ݺ���3� �*���wz��Vֶ�J��+|5�Pҷ��+a6}�[mZ� K��(�~v���Y4i6E����pͪ���]��Wy�JK9T|'Яf��*��`��l�E��ւ����ǂ
�S��h�T�i�e��N�E�V��������M����������2�W�_�C���`k�~o�m��}L��|�ҘZv*b��QGJO۲�����}-����OF�<��̐�E���8��@m�F����e����g�U��D`H�Ŧx۵#������,52��P����Tr������t,���~@6Z��q�ސ�{�Q^N��G���ȉ5���K�'�Q1�L3��Hň��2v�A>�e�����dH(���L�g&�a!�ï��B��H�f[���� ��9bvh�q�����]���%�0/d�ܞ�k�Ɣ�%�"�y����l$x�PG�RK�.� 9>�4��e���u���/c�/�D$�	0{lĄ�H�8�)���s��"�~O4�N)�f:�'n�-�E�=��F��� ��e��Q�۳c@K������R���x`f��f�47��hܻ���4	Z�P���I�VO�y�n���^��q�∙@�	+�&�ñ����nE�ڐ�5��㿛�|�~�w�b�c���N��3z�XL`���7�҂��+�8'�BQʧ��	�2J2w�]��{D�`\T��Ծ��1Bb���-/௑��g��v�Tr��g)�b�Ȁ ]}|U���)��	ȴ��.V����J��$Z���`�y�8�;�7�S�# 4.��³�f}oH�^:�ԏ-��\2���>���%yi	1��4������tx�
��HK�!L �M:��J;]��^�W ��/J���;�i��(Q�X%���� j �*���_��|Ck yV2�~�%����"��]P�����~l�-�l���_�Йg�&\���)��\}O|��7�n�Q�L)��fۉ>�x�!}��n�d�/�z-F;*K�O�*7�j<z���M5��6�}��3��AD�h��C�#
�pE����^ (<�����#i~�?6W��*��F�|W�۹�X��K�[�G��tKbZ8hY�3�,�H�=��ܧ�Ƌ���a 4h���[��5��?j�o�T̻��ȱ�����K���#�-j��^�Z�+�؊z`�~a���8�o��q%�iTG9:5oo���Z��Y<fl
%`�������\}��Z�Q��͉��V� O���Dz��|D[�Q�5c�+��l���{����ga��HX�����S��\���N��Q���x\�,��r.��=�,;�B���'�o�Ƀ��⋚�P��Îd\��ƶ��_��2>�K��9��F���
��Je��f+%@���!j]U���1�	���E���)Tݻ�X+{�Y����{�@8�q��K��Q�n˒���os���-XjT�(��)�:!z[]�m���C,���h~�%�ۆ�V1@����;F�l$�p�g��l&yr��8G�����9�FA�{+�g�rp�at�(`9i������A�u}jn�GI	#a��":�S����vL�����a<�����D�8)*�I݀�?+�����>,���㜈�T{��k|��<J��Cu������/7&\T�S�J0`9d��Q�fO�&�:ۡp�G�7��"����4��c[
��5Hf�Z�0��Ө�M5K��Ts�Sy$*���>���J05C�Ll ���T��(�C��>0i�l�W��;�A����m�����T׿��۞j�s:@�d���hl����1���S'כ h����Κ��Ɉ�[���bh <A'���Y,�6�Z�zÂ��@�TQ�f#�%G�R�9�Ǖb!�������a6�U�;4�J�� "u*(��|%	�D �B5���eJ]��}��U�i��k�����x9Q��w�kʔ���A�2�^�V;JR�a
�;��#2vǲH}�ʳ�Eq)��k�W���D���ܞ~\��x�ۡ�����B�8�*j�4�pz��>V�h��M޿��m8�B�8Tɷ�����_���;���+��}C���Õ_����6��d�"tkK���l�i¯��U�s��#	g��t�Xs��`���Z����zA|��� �JR����F�4+�o.d��v���u糁ć��i��o��uM��u0�~���X�?T:�C��M2��U��/�;y�-=�Qq��2Z&�ܾxT׼A�b �[/��_��`�q�T�4Wۉ��0����H���h�w�O±�f�p7N$��Mq�"�x�&P����f�}Uп���1�cg̶ ��@��K��k�pH0��Qa����V�;�H�;oي��?��O\r~+J YrGWB���Z��$��3��ML8s՗���*rd�à6���D�b�Gϔ#�*)�y�t w�WSquYM담����{�zR��ߏ� �)�2W+ojǳ��L��_��>o�G���@(ԹU�g�٘�'�O�Y����z��,|�s[�'����{��*���dҫ�UX�����cq�c��S�/N�W�;�C�c�_A4�CԟC,Bmn�/���q<,���Z��t�6՚�K���}7an�)x�RI7]ϒSʰ��&~�uz]k��;��B��4h�<׭�u�;��>�L�ȟ�K��]TAٗ!8���mf���R�0q}�7Q��Ƀs�r]n�%9��"�`r�?�D��qw��=l���y��4�oN�b:Tn�p���=�E������#��oo/���n2�����_���O��>t�:&л'4�w����9]���i���z��s{��4�������mKq�C�1/]�V>UD#t�
�ϨX�i�.�/3.�S�H�9����pC�	��e�+��\8QyY꫁z�cr��gCւO8,+��E�����9>�<�~W��'UӼ{*F�W'2����EN&����!��W�VG�������3tz�_P���zNе+��~!�evi�o@O��Ɉ^���k#.�2xOOU��t�-I�s�G~�_�������d��n4 � }4ѫF:f{�4?0u�c�8ޢ�|��~������&�m���#�ퟓ�ު(^U�)��L� ���3~U!�������ҿ.43#8~Mٶ�Y[I\���&Fk�ɔ�[{ɍ$N���J:��6�_S6�EŚZ&W�Zp�g\�������;�?4�D4�.�gv�k�l���������BV-���4F۲�<Y�W}jѡrۓE�;��/�sޠ9�#�����;JM��/(n		D�#.���准��}ލu�RS�ۏs��ccD��@�i\���%���~��Mx�$���ĕ��&=��O�G_-^`�4�u��L�K�"3��o�8|��M.
u�b^���wTs=��Q�n��-"����Y�era�@Y���lo�sr�P �{��4�˻VĨN+��VBq%���4OI��j�.�6jZ+'��=�\_�i4`JLs��/I��-(�K9��u�I55D���ߖH@���4��u?(Ղ ?��'���-ͅQ�{�-u3���vc �v5�N��(b�h����lα{W:id�Ъ�	�O��\2���uL}:$��G(��kz����?�E��'�#�h�F�:���i#`%��Mr��P���d��J�ƞY�m:��>p�W�{�������~�D����.�@CZ�6����=�,�:��u)Qw;���χ��ji[aꊿ������|��'����r����V}&y��~nx�4�<��+|}�4gѶ���n����ȁ"橯�:�
ǡ��I���H�bq�ڲ{�7^��?���<Y�F7�=�Ҙ�� M����������ec�qR��f��NZ��6���x������#�q�����U���>�u�l^�����<�~ZI��]$����r��fh	1I�����?�M�{�$ע���ę.�^ ��}�ؤX������},|ل� ۽���9���Z�i�8D�������\��f2�����;P0�3&V<F�y���tU'f�p��;��)�4�2	
=yAѓ���lV��x������:N/��&��+��z�דC�������?k�@��Ukɬ�d4�h̬�T�Wk�3?Uht��%RY���F����l
V�D5�����J�JN�I�Ʉ��#鍔��S��+�#9�mgƕ�����J�O|z���V�o�!�\")*�W�G�G��J���j6�LH�G��zp�7���!Ѳ~��*��(ᢥd�_,����Eys��v��r��>���
���^��ƬN6fq�Yj�*~��ʳJ/�`s��O�ž����g���gY���i'���d�#���� Ac���[¡d��_��5���<jY��X��V��������p�z��f}��+ݹ���;.5�/�� ާ�o2y���;�-i�40��0_<�؛oİ`8�H��5�2�k�X��V���p�b��NB+H��,Is�=�0���B�r�wG�OE=U�m>r��a'��1�)/���&��zWCwF)�gZkF�d�����ב� �ƅ�����}��(,9䇻����P��W�^�ٻ���Q���IQA"�Ԕ��s6@䗍}�@����P���Na��%3��C��=:�Wtӗ%Q��Lk��YZ��	!\��r]���G �2��U�G	q� �
��<��H� ��l&��!��80�V,&	duG��j�)EB���/w���_F�ौF���sFai��,��P-$}�/��r��+�v�O���s�h�$0��7�����M�ÝUb�k;_C��HT�T�3Ph���-_�&�O`�~���A��bE��"Ua)F �6&��Ui�JDmUR�:���g��'�w���J5�,E�ō0�|�*`>��}jm#�g���� ���RP���iyp�p篴�6ީ)	���t�Ik��3NA�;���}F獳w��m
�������"FE���`����ק=�>�M�{��N���}WA%�w+I�䃠��?BxG�s3�X���S�
T\=L�7a��J��k��Ra�+L�����|v��Kb\�jGp�1��i��J��Q>P>��������W5�����7��w'��@�jƃ���|�w�n�q�?��%�&��ixC7�4@�Z6�/C;��%�+4�΁�����!���*M:��s������r��Z
�P�"s�6��]S�G;ª��T�H4��l/���s���
���y�/���hǛa����,�:�x�����]�ў���ip���v�y��o�=1{�R#�D���r��g�'��~*��|���7��ʤ�t l��qKmiZQ2�Uuv9�����άBJ�V��͔��m7[��
6�(�%6�ɞ}��H?�C�����}����� �a��ɬ�����"� [P��%��%9���0r6[��#���ms�����i��kf79��LS����A!#�q.z�j��3<�0�c�N�+1��e�F���Q�m@�)dLeGm_���;N�v#��S5�J��ԐѪ��:K���~r�mSp��"�f���W_}	|	Ճ�p��"|k6��PI�E���F�+e@A��m2W��G<nf"y�'� R`��][�B��.��
+��.��|��J��4������r�?��8�L���"�_;�U��O��xt�	G��wL7��zڿ�w6�5w��(q��sf�ɨ�c�l��\�z��Pv��ا�l��g�T�6KL�W�&��cNn�.�w��t���$�N�i-T�Q*L9��2)���
��c��j�Q��Z���7 ��?jW��QI�d��:�ZsP,ky�(�U��V%"~�}�U���R�Vx0��v4G-�
�[��-����G�D�q�fVc����@{8����dz=����N,f�<S��%Ϩv	#�^�.���sG�m����;��%]�z��w��~X��	Y�7��������3��uNszο����-n��4�8'ld6Ecq�ά�ڠ��|:q"yuRn�������\�V������9����H/��i���}��6E0���B�y��E.� ��������EX@ФDc��梊����xg��h��9"������V����%c5��-��~>}і��)��c��?�c��˿!��]ÈXw���$.��S_~�
r-<�jPН|�K��g#�����2a�o�,_�����{�1������*�B �'��ޭ�� �#-Qey��#�l�ӫɡ�L�����l�}z��d���O'�Rf�l~{i�H)|��<Ht���gO$E/zrn�Rh���+s\����Y���ˈ2������91k�� �t�7�Nt.�/¿a^[���N���}E�b�=L�D�^r-�����R�J�躭� ���i�������>o�I���b�N�.W�,��b��_���Z��l���b��o��{]�jr�\F��YG�W��x�^5A���Z?��\O�s������O�Zsa�	���e�l��٦,r��g|��[���k�׽Z�כ X������%{�
�8�/w\,�?�O��I���� �P�3/��4�����6e2���U�j�1]Ђx�_��+�J�����n��Ȩ�Ղ�u<O��r�Iz$ӧ*k5 ��#�tkk������\TXe�����F�$���M[���N�@�}�;�����iB�E�1�=�d��p���iw�d�ǟ������@�ljT�it��;�;�=�w��^�}	�[��C���uF'�"����a��6Rׇ�ΥI̸%��.2��� D��)7z�������~�������+���C���1пCe�"/���{b����x����+8"�!t[_C�< ��mq(�kp�o�X j$�V��~��m4tKsq�3���3w��v,��x����Ӛ��N�q������-�f)���"���?��S��y�DCa�O��mc����W�^uMi��(�.�n���]wh�����<,��v���ּ�3�>�m^�os��l4�2��t��_^ZQ��N��Η� P�W��}_��M�_ {��k=.l���L1�/Ql�*����
���leyi§4L}���\�p}1_ &e�,kjV&o��1�-�}�$.N� )[��!����]L�3f������X����"z϶��a��i�d�~��+�A,�ic,5�K��E�麤F�O�:�x���{s��络g�׍��EB3T5V`�R+��MsMom/X�׳,�?S&�+��t��1��q=�6�>uL�]�)%H��n�I���I��s���.�GJ��B�LN�	v[�a��粽'�pD�{��<[`��At'��3�$��V�����C��P�}�&r�W���Cم���p�@h�E�u�B���O��|�Ɨf��ԡ���ͨ����T����i��������kvat}���G�f]3K|ƭ���U��u�:�u\��o�;T����bI�Uwǹ�;�-�^�&�mD1�ݓ��a����	�7�WA�'�_s��L����A��@�XX��h}��=��`�m1����狅�!��h8'���_����1�6�D��g�4	0�A3AA&�ʂ��e1m��:�I�u�?��O�H9��!�ء��鉋�f��(+�⊯f�w�d��ixT��)��4q�(����(4���ҒC��zp͉�D��K��0�j����Īh6:�V�ᕠ���X�aq~b��C�<����ݗ��#��Zu�hƻ*�Xa5��%����BY�s> �]���#�Wy����6��|;���y4t�#��j)�S(G]�Q2��Fc��}��������1r.�f>��H��P\)aJ���gA0�Y����h�`���@Fʇ�V!{�+;��c��-씍����
���RL�P�	!A<:6�u�v�����b�Z��^Ƥ��"��ͣ#�p_�,ǧ'��ě/\=��c+UO3�m4폥zsbxE#n��zB�^TO#vyӊ�I5�ϡB�?�AVY�v�1�(����yhќ��>[���@�^��y��vCq]��=]�U2�ͬT�5�'( �]j/|����m��*����J(���fԇ�4�2�Xa�jˈ�/\G��خ��Bt/׹�C9L��n?+hdK��8�5�e���+��(ـ��7��b8��JS�	�	���j��̭l�x��d�PX��fw�r�ئ>��>w�_�� `6�?_��9=�h�f�Ϩ��P�~�s���\�c�fL�0�t�m~5��p>�oֵ�7�����7%���r-)!�j����&�KO{C�^Th[��x{�OH�N�I�eN���ML�9����[Ț3Ѱ��d��_����eq��X�����M�m�S!�YWV��Dd��<K�v�3�(�v��"١n/��6n@}���N7�f;��$�Z�k
o�z��I9<��̣${�_wt��-Lݢ���v*^�t�[��k�Y��p�ќc%�@5�
�m��=WQ~��\�T��ê��7�N�y��ڋ@���{�mC]5Q7��+�}�$e|5����dG�ە�;/�f��c��@f�:�^w
�#;�P�"�*�YS-(��m���{U�Wp�ƾ>w�`R��K��ϽG���dV�A1˶K�;��<�g�m��R͟��9�K�#��&l����,�}�u�����D��M��ۡ!��h�[V�U5���q�L����i�a>+1��
3a�%V�g�p=|��:@�鞲���ʥ�ʿ�è|}�F��@S�(�ă�#�?�r��bK�����c��������E�MQ9�-n5��:_���`Tf�k��
nX���g���V��*�>s�{b��:��)/6�|��-��,�%��/�Zls=�R=p��z]"�*�P��wԝ̶z�h����х�l}�
V����;L�[��	��o�C�#\.1�U_��9�a�,�,�P翣�+82)F�]DU�?�	����m@�
�����D�����u=g�GK�e�eq0���j�Bq@J���������U�}x�2�}�]���SWy ��^o>C_�m���jUU�^�_�Y��N���&���
q�0���ݣ�Ɇ��[/@�aH�J�J��I:{Ѯ��I�tWs?����S��u�$N��
@����}�L�����Y�h��m#>���rz��_6.�n�}z~�څ0ͷb�d_y�M��ڝ헯4jrV�ѥ|� _eoDI��p��G2��Y�Xq.a�����_�b��,�#�7��:���ׯ�#�E�P ZV�5��G��ݱ����Y�Mk)J�@{����x��/b9��6VE
]��`��k3Rf��0����_]�u!G��"��bd�R�m9b�z�'V,��@_m �@~/3r�y�/�V�<�[��ب#�)s���]m
b{rM1���]k^mV�Wެ���y�Z�g����ԋů*�W��5��]��=v��hs����|��}��@O1�f?Ú�UQ۹��l��|�yg�g@mɅ���fU�)�	=-�)p`z���Ϗ���<�wW�Ǥ��}%~�w���� "H�� ٟҞz��,�s���WK*������Z�M���$X�NLP=��[b�A���x�\;��#$�t�Zio��d�.x2Ά�7����~�@
^�Ny�w�Ms�MTNd�i���)����.a�l�FDi2�4v�o��.p�)�����oX. � "������9wzȍ�K$��C�)����	û����O_�q ��).�S]�n;+C٢��Ƭ�"7��] D��ؿ�Zt�D����:��4OK3�����t�?��R���H�-��J��{��0��|�-��M�MۚW�d��&Řj�wi����C�O5��W�a��w^�
j2�[�t���ʸ�p93�����C>�S�*���ު\�K���f�s���uE�)9㹠���#ʏ$! '���=C�,��ij��&Љ{=�>��OX�J�IZɺ�� K��S�[�ы�n�ϱ�OM��e5f>k�M�8a�؃���>�0��sHj)�W����"V*�)��e���o2'�!�t�<tY�?��JoZ������Bٍߟ	��Bѿb�N����H�ˁ͸����%ba҆R���h���YLXh�Gg�6��`	-,t`���E��q�߮��˦RNVO�=�J�2Y*DɊ��T�7.�g��9��(��\��v�qs� �������p��e�Q�!Z�|B�B��H��ш]4Z&88a�Y1���Hp�O��ʑ{��W7������G��$o'u�䙙9�RϏ�u�H1M��/�����f��L�dF'E��R�%JI�s�?��O(H�{R��Fu�F] �b'qj(=�q?9"h��#>�$hfR�<~(�LY�a�!�����.zT�JPْ��xgP|�Syӯ��i¦��[~@�h�LC'b_��*��m����u .8�<�|�����r��K�S7l�s^.E�.8���*�F�yk7�M�%Kw����M�K��J��\YU?/{��2���bQ�@qȇ��^^O�Z��7>����� <Z��E��l!�(�s�~� �9��x/f	���1·��dO���ٞ6I���bNKn�Rn��V�����H#3��F:����N*��Fþ�Je�
~������H�]��El�����}k��]Z��Q�1g� bT�f��{4B�ZJ]����� uuuG�D�g��
�c6�V�#0?�1��Ot>v�L��mPњUe8�V�)?�p8fy��X�o.�6�+�5P�����ܧ~p��¯3ӕ�*&����F�mD�{^����/������+��j�жί�_���]�(_���T����WC<��)L�]�M�#�	�X���p� 0�3�s0ײt&��ts�2�sf<!���WS1�����D�j�y���;Q��B:��@���������9�t]�c�8]�)Kh�ǹ�x}G���e��#����� I���'�Y���[VʪP,��y�i/�|)�^�ZW�c�<��7�+m ���--���c�/�tĨ����"�^Ej���f��A���0!� !9 �Z���:bǤ:�9����^���+xT�|��w����9.%�K<����q]�8xs`v���9��g�Pk��A+>�4 x	AK�Ft\"��Kt�8ca#�o��{�@E���Ƶ�Fʃ��I��H��
@{�vK��v�H�4�p\�r]�TkVM6�^4'P��.��*��HL�hyx�����I����bG,���>����~� �JE��YAs ����2cF�A�ݓYٽ_�>l�t�Kw6ݽU��2	S�j��	�6�f�dЯ�#M����~uG��@�)Y���q`�w�Z����x
�e�&�yb�m c>�\N����s�ΚJ!.o�_z��Ǵ�ʀ�kِa r�����-~l4��7����m�&VC��5��yt��Ր��F�|���@�V�y�������x{˰(��}EAA)E��a(�a蔔ΡS��Rj��Z�%$����3��}�׹��s_�xv��ֽ��E�?�xT�� i�-�ӈ����m�M����G.���hN�����?G�����Dx�q[X��eY�� F0�9�?I��Q��T���?�!��t`�^w	Zq)۱#���@��l�LD��k�h�j���=,WQh�G>���rr-� �o����`/q4l���S�m�)��ϒ��*J��I�,��b����
�$5�Z�-l8���ù���K��t��n��tz��us�.O~ ��g\�l�j.43+�r��Q'�'��j��!��̡c��Fi��OB0µ;Re ���L��c��ݱ�D�J	 ����լ��D��y��K��È=�k�I]�)��[�AcW�˰��@=;��Ф�l8lhCO�ZO՜'�0b��p����xMf�=�)~�m���f�k�ԏ��Ma9��%�D$1ܝW{թ�����"+�k	��J}%�>�	�U��w�C��<wT����.��'6u��f��ؓ�<�����(��@"እЩ�n�c=����n%�>�� ����Ck��,`Ҫ����5��A�B-}�e��S�:��[�@������j�e�{b`����ҹ&�_���*���&�{lw�\�w�x���\c2�#����mE�����Te���]$�����Ef��7����2;���Z8�6�O���u�ב�bn?�x����7�[�$G��@?�eី�B8)C>�ɏ%��B���J�Y�+��˄xZ�7z)��Zit�z@��`��]m�����eZ���UT�h���z���8�oaU��R�.L�_6X1�ءR���>$��,�LH���{u)Q�����~�6��p�1���L<��B�,�����q�m���;2�#�ܠ�L<��֝#����c� �W�Gs�2¯�%M*;��?�%��`�����q�cF��� |�s��LĊ�0�M�f��^����ma���4�p�/��������c�k�A�=}M�M���4%�Ut��8��g\��62-D��=띬2��cW�}�%G�	t�핁o�Ƅ�Tb����K���@1��	#U��4��K_�Ej�i�����F�t�n��J]�e��-K>�{Fvr���n+�EW#�����'��[q�{�H�^N{_�d��p�mw�)�2�O���y��h����͊.��H��z�αD����#N5�������uk�\c������<1HG0�2t���j���绹w��jUkV��!����Ȗ��Ǎ�l�f_]�8�t-�wP�:)={��)*cF��5��|�d��
�2{�l^r�.�~�����[$�X����[΍�%�	R�h��ؾ��gp��Dw�����|�:�e�~�$_�,�T%��S�-q�|�ր��k���0~����+����l�Gp۲�mN&ڨ��Ww�f�>�%���غ��[�����X|�F6o_M16��_w��]�֨U	_M���ŝ_��0ԾQ@�r���zڍ�����\�?�Pym��~ya��Aҝ��P�X�[�(Z���Mir�*� ��krڹdɫVv��s��l�j�|�jx��Ɉ {/p4Q'B�� ���Z[����X8�������Cq�<���2��`��8��ӝ���\���t��jp̆�F�N�t��V�oS�w庚6�#���n��� j �9�V��@�v�����\�)����u����c�K��`��1������� �Qbk�kw�K���L�C��Й�g�+,y^KM�=խ;��hv뻲���������ވe_㭸aP��{�q`��̴��'p[ȴ�/�����_�@�ݺ�B����=^�%�5�Ib)��6b}O/3��m�]��i_�_0�ꯩ9�l����rן�4�cZPu�^��()݉���P�����7T�MWC��Ma�24Q�=%a���1:���%��%&������ǇѢ��)b+����"e��V�T�UEw�r&��̅"�̅rˬ�����m
�G;�����| UD����ݞ����1gm���Y�u��z=��]���ɺ�?]X�řŞ�Po�tϗ�_Ity"M��`3p������ń�k��P�%%4��C���U˛%8��c�'�q�B��#�Bϟd��1=���3�|����ki+fv󯩂ه�ܳ$R�XS�U�׻�8ÿ��Y�%L����#G� �p�Ь[\W�(���PX�u����.O��Xtq���As��:D�%�X��xqAf�"L#�f��\�0�2?�j�+���#v��"z)��i�a�n�"-�Q�	��K�{�4O�e��!�ı6�"�S��Z���� �:�^��j��t�ݪ�u	�_6��mw�K���F�%N`jD��"wgF�.U8�3՜��q�"(\�6p�d\�Y�&7'��eGkk�no��wL�|�y4�o�TÁ���T�ހ���F`�Ը''-P�>��)�b��������~���#�#���Ѣ��+ء/�gOsR�Z;�;�>V�i�d�N�2��zzj�f�:H˂z�ޘ�JcV�M�-���=�����l�scrY�|9�`끫p.(w��~��m���FNQh�.��JK<�Ko��@	�pKo�M���3�$����Q֚�,n᎔�kB�k��O����l���n�5�7o$ f�.��I�ý@]�HZ����j����<(�c�F�`s�<I��qT�(]�g������D��U��X������KƝ.�)N9@���]e;��殲3��Ә��# L@D3���������.V�l�	n&F���`�����|��2��J�R��C�E>���������y�Qc4��T�(爞�����{���M}:�<��5nCJ�4�ɖ���;�T�ڵ�f���vǲKM�H�7���ܬ&��RY�t{�S������n�UOx���SV7��8I�+h]{�zf'r���~���t+L/����! �3)m�zº-	<n��:=���#�����4r�>�/���8)'�jf鵤�*�VN�=L�c�+��g�<�&az�/Mvd��[�S{*S/�P'H3" �9�6ꢂ�����I��Z���֗���������[�H�n�Ƭw��ץ�	K��Y���9 -p����^.�P�ܿ�d�3]-sA�)V������h]�o(+S�}oR�X���G� �Ze����x��D���BL�N~�	��6�
� ����Oz���^�����#N)�N0{�|�>)GóQ�s�h�8������b���B��_X.0=YΈ�[��+q0�L���A�](#n���s>��(�K�����}�����y^z��	~h����Ot8O����u����qȗH�V������̉��)��+�Z���A[�--z7P<�=�7/�mS�!xE,��9�E*զf�<����1���e���%��n�|c�~�,>e���~)����hP�o�7�nF2H�7�qQC=�'�����i��2w��,]��"���(�\�����_�@�?x��C��c�N�sʸ}_K�ldY���(���>x`�[z_���a/��7���<$2��^���1Z+�:z�!�M���߄_���h�����tTY梉p����8TҀ(Ш"��5�������z�NL�L���y��X��{D�F\�&.Jjy3��{~�z��N&�V��FfW��=r��Dvp�(G%��hn��ux�oa��~~X���A�,4�;�f��(�'�",�܃vr�:x��1靮��1�$�4#�¯f�#�y�������:���c)���4�^��w�l}�g5�����8�p:o���9vҲ�"�P���0�u.d�;�s��Z�ٺM�#U�1�� �8��q�0�03J��u���Gz�r/��J[�o�V)�-p�wN��9�#�	�J�� �7	���|
�;'a�G;�qq��S��
�zŐ��2��^�����H��?%��+�m7Y��1�i���T�m��O���7ً��nU�[H�r۸�*%$7�t����m7m��NU}(�0C||���n�#�5V�؂�� �
\��e�c�A���X��g�W��ms�gyJ�` �gU%���P?���L��S�j�h�!4�����T9�<�s?^���z*us��iT��n)X]]VF&�p;*��L!Ftt����O^��qn��i.R�H��&-8�������Z�B��Ɖ�[3�%ǐ��g�&�>��l
mRZ������ZU���F��(!�1�t�4n��p����)�DE�}������u?D����=��۬=����<�Q��u=u�6B�-�堙݁��L+�d!�~
����V�A���Z�#>ZG�>PMev�H�q����YIR >v�(�}R�"�]'yw��'�=7]8޾�X)�����2���8p�A$N���/�<�	Uh���1�j\SOb�c��.�Ǝ�e/�	�h3T�\[[�-`�G���$_?�-�����de�¬d�L���͙_d�	 `��� P���!T��{))zJ"Y--�B�7¶�&�����8�2C�*�L�X#K:n�[*+�Ľ�o���ּ]E�~,�	�û�Z
ו�~r"e��f~��(�)@�;}��@�����v�@�Iq?cP,�K�c�=���đ��8��9F/Y[�{�0[��4*KkhT�����d�������_�ѿ45����V"
f�@ހ�	z�sV���ĝ��
�������ك��0���bN�J��M�_�ۤOݖO��,�GHCn7��������1����&�4(r>AP"�o.�rV�1K����<�{x�fk���ʀ��4�I����޹�L��+K:����,�q�!av�ϛ�8~�3������K?k�8��s�E$�ˣ�^����#?D�<籪T��U*�*��E���U�Co+���x��Z`e$��C֊��D�'���w��.���Ȋ�`����:�c�/�zڞ�;+�)��y���LHe������aOR���90������|m_C5@F�Ÿڝ�~�E�s�[x�s�DU���*�������P�v��N���*��.���b�B�36g�E�d�	��M"M�&��7�����b\�/s�:�2d`�ޯ����'�dxۥ< �����fXCPppny����,x���0�%yE�N7�9���0ڏzD�Cuʠ�KKK�'�YY�q�n�$<�π۔� |���Em�xq���ҵ�!�����,��qq�^�a
.7���ᑑ��)��˹��<�~~Ɗ�
L&��ybG�'�r D�і��j\e���yyyiЀO"��) �f����|^����ͳ� |�l#� y%%9j5��B�`��� f��e����`���{L�����n�L 2 ����e����������M)�£���vCC��o�}�~I�����&��vJL�-}�p> &�?�8ʖ�*q�����q�e������V���M=��Ϸ�D����&���	gr��|�����~8�����f5��߫��_��jaB��s���[������l�.�u��f�[�JV���IH�Tۉ�QB��!�������:���<'�e������<����+Q������QC�}���ߚ	���x-�?��.�E�~k�~�Qzj%.n�9��T
�P�eQ�l�O~��]��B|�]�K�b�r"�SeoE>�uM�tVX��2@ǟ�I�(y����2���7�(��C8���8y$���h�|e$��8%xFɶv}��������P���Wf���^��Z�
��W�'/��j��}���N��a[��&�A�S(��::���L���~�KvN^�P�&�,�뭝.�����%�%�yHy��߭I�K��s�.Z�Y�d��� 3x��>���*�bJE��T�} �έvZ���I��!�m#<��\��;�$ϊ��t�T��*h��vY��H��q6���z@��U��w�-�,���{O�D�@�l�~���lą��;�:3��n4}§�%�[��Y�ټ�\kf{unꄑ�?�)D�d�f� �����f��g�h�;��"�3c��ҡ������p�e��{��[-q�����b�#��Sr�X\��j &������������\.U=���. ����SE�5/�( ��C���*�!�h�kL�>{ >�C���4�#1��q�s��� cn��
�D^ze���]� ^�jbY�7��>iU��N;>��Njq�q�=�Ű��jsYt}W��Wd`��H�&��xY;�D��瞙��z=weg�f�v��kWQ�a�y��ф5�k���"�ئj���s����P�ꏼ7J�h�q�O��'�sZ�)�
���e�-�y��JS�E�o�.�2@��ž�ҳ��������{��Bt�]J��X}\~?�7[X4�0W:���׺�r�'jSg���8�r7�r�&��0uH�e-��D������O��?��ƺ����N]��S�� f�f�-�4�D�,M��':A���a�������aL��}��o�I`ht�#�5./��%y+���	�z⋲�S��%wn��Cz�x#!"�Y�/�׵'^�#��f?j5x��
9F�H��R
���j9]�$��W�����I�!̨>>7�'pW؁�{l#���@��e�P��⻸'7��L�F*b�
���,�;A�K�d=�i��[����#÷: E�h��*�?DS�F��X�5Uk3z��JR�Vz�eZp�Rg�T�}BJ�N�A��]qX��-W��tx��&%���RՉ����#�Fa93�H��2z�kq���j�E�gX"ΥH�?�5��?�Y�_�sQ�*ވ�و�˫�m)��:���يXP����4��d��Ok�^���^���4k��_oD�Ǟ��cr=��ӝ�����7
v1@@�1�������
+Nz�ӭ���nw�f���Iϱ�V5�O���c��;U�i���v�OG"��m�= �x�����
G��ѫ��.�*2�h�q#���/��G�������嬊���_<��r�'|be#e����a�y����ߩf)���!�C���&�OG�yȠL����ua�z���C:�U��"���S&3�=�6)o�U�8��k�������F�R	�z��k�V>l��� \8�t��7��6
�|�����0*�����`2���N��;�{#!�^�y%�o��:�-�����c\dr��m ����3k�i7_=<�\� ��߁��2���λ�Z�7�L~\N�3.�������d}���V��]Af�WM�F��oQ�U[�d��~s��s'v�>�q3��U�w��>�y�b٭c����&��Ӛ��#u����y��C?�b�I*�W����M����7�B^�Ό�/A�fu�=y�	��3ls��9�B�<^c][�wC�`���ѻ��!`+Y�5����`�qj�G�o��6<��~���FOGJN�b&�k'�oŕ�$��C�}�?*�}D���R�VN�@�*CIZ��B�D�����2�����Q��7�?�Ey�VK���!�Ce�yt��~g]�ie�;�!-��t�<1���s|�t�D�A0)��_�h�����{&:<��E$�%�J"�B�`'t�%F{�M�/q��5o�Đ�s̹ Ю�szc�s2��09��"�d����v��!Iۉ���@��Ϩ<֘hIV.Qm��
��*���Ze�!U��R
�k"-{��g���I��x���6����r_�������g���Au^y�Ĭ@��
��$i�դ{\���M�*�0& � ����WOsP��[�1 pNB�����)���JL�DIF�.QD|���o��򲈍��=$��
YoK�D-�t+��>�F������&�|=�HlfI�[�=��I��5��Vk%�0���K� �X.�L�����RJYK�8C��@���c]����#���ز�o�mGU���|�������p]/H0��<���=�J-�[��'����^�x���K�O}�7M��N���R���g)Ԧ0�|P�4�{G�C��%��� h��������|��d	W�=^�`�I�h&*� �Zм.GosZ�b�;<�VZ���GOI��Ӷ�z.E|F2��N�3c�o���p�=�ur�!��;�f��2ae2.E���Fy��x���I��9���c
ܶ�f*΍/����b�K�}3����s4�W�Ne�?��p:���A��k]�kS'��+����`���.��$L*��'�h�t͵�Ԃ�^���/&!}�C.�{���YҲ�S��9��a�p�]>٬*�#D�UI��7G;db{xr�	�rI���γ�n�"��`G6g�b�pa�S
|&�$���߼�H\�=� �v�3��F�j����L��9U��(�K�*9a�:��dg���$�:Y��;���]$d,��BK|��6�h8Q���.�A���ҍ;g+-h<$�@{4g�H�������Y��\����l:Y4*��l2E�g���bȵ�y�l��k�h8�3]�-	ㆴW��\Rn
�p�����@Ob�/�O�ޜ�z-��zE�]�(!$�i��m����2^"ԇz�X��:�چe�u�זc�Au^���U%k�jSJd�]��Uõ� �vR_G^�1!�Yt����S���k'�?��Ecm��vȊ�TUHh�-����!�WGT
@m�y�y7G�Kt�P�v�kk����N�z�}ݑUÎ��j���-�����ɷ���R/N�af��7��4��7~X^������b���V�X���%&��@�����a��q��i��P��;L_5�
�<��kR���mՇ��B4��݈@F9�l~]��˓B�����zU�m/t�����Y#���P�P.�S��"��XJ��MA���Z���-�Y]�+���r��v���9�幌�����"�zN�Uc�ka�TĦ�if�ߔF����Š�D���UH�V��Lv��aB�]C�~�Vp��깯ǀ��S�)�}WaH{��ǣ��T�!�R���m��'����O���.��Ն<x�2L�s}��qZ!
ځ䎰�Ud�[B���X��8�����X�3��W�(��ۺ3�֮75[�?�-\�0ˆoH
<��bm2n9J���ƛ��l���95�f�О��_hUY�������'�9JS�*@tق&�B���6^�BHٖ6��Gf8��N�|���lR��#�t���~��5�ƪT�O�l�����]x|���J8�u�C%�@���#���o�Vl�dVmW�	q֔��HYE|�&��3)5a��ВjWC�d�+��^Li�J�(���iׅ�o�Ʉ�����84y���<�G�[�Ch K#���G&<Y`�S*��G).�G񧪏|g�2 �%<�z����cX)�r�kP�;x����H�?d�|��j_?���k�b뉾����"�4mF��aW�U1��Zx�9��&��c'�� ������i}�{�٪�3(~�B<)SͿ��?�m4P�|�d������JIk���莇�R[Skn|[�(\g�������
���1ڤ?������"p�c��s��4�('�*��=Y���s�S�l�*p���zT���~.�˝��O<;-	�>9�Q��W,�-C���5�G�f5=���u�14�A䥇�m{`�۾F�#4�,}�tD('kC�9�cP�������g������
C��5�?ς�Ӵƹ�˽�U|�<z�5�Љ�jC����
�X)���N��T�T��G���ZKH���M=��Ͽ�\.L�Z+G(5�*�<5��|�F�u�ŸϺ���e������NE�Z?(���N�@B:������_��Y"�,Cn��r%8b{�y'<6�����$�<ţ�=��,/�Uyz.z��*ݭW��w�!v�����kX�\iK� eR���<���n��t��1Ԝ���+�1����e�OQZ$§�魏�P�mב�Վ���	0�~�Ȧ(��d�d�����7�(�j�G�'�W�����'�T��l����[;�Z~�\�����Az �=y>g}��.�W*���ć�q���>L�;Z�(�V^��~z�q6ۃ�Y�|�T���%�]Gj+Ou=��ފ��#�	��#�L*9;ע��E��E�~:���'�m9��I�%���V.�pܴ6��VA}��HT�DO������Ӈx�`����)u���b0*3��L���d�x>5���Z���,��O�ު,�`�$t�H�{=�Dy������-�_F$�:o�(�t�P�x�IB2a�G�ݙ.޲�ڝ�2�*���\D����%��Xx������Ad���G"��v>ߎ��Q�v)�P�Wl�W|�1�� >X��H/�����*�~uk�p"QAj�9�pI.t�o�����Pťn��z�"D�7������&�ԇ�Rj�Ϡ��&��A��G�4L����	�[���50�{0�WLQ��?�f�i=OhL��殯y�6f�꧲P��U�eٔƺ�{���:��I��	�ߔ{1x�+��&�6|����G�ʪ��S�Ո������=t�BF��g;�]tp����Y���s�o�����9��"���A蝜�s��lE��@�Eu�;=��� ���?m^.B�[̻Cc'�5�"���x�@D���㉘���Gq����B-�"&�+�h�l���z?X��6� N��]э<��%�40�l���
!&���;ಹ��%n�������I�~%�]'Q�׵:��WO4��8��ym�+�l��z�7��ڳc���q=������j��z=�A�J#�v/��S����3�@��	Oڍ��w9�0�Q��Q���>ѽ��4+��f.rw|���f�(�;۹$IV���ò���Vb�*_WQQI��̣����g��3r,e�B��a�ʷ���]�Y�E��7���ET�' ��"8�g�l��_ow���B��Hmsm;�`�Z��^���ɼϘ�j�������u��K���0�މ�HF�:!�����?QOI�Ը�O
��]e��/�2�׵��\o�;�SA=���{��g'���J��|�L6�w'�vz��5��A�T��5~'Wk�Y2)�W�3$�4$d����zτ�?j��;B��F��m�"���y�����k�تX&uwk�7��j����ދs����^����A"د�|�؝TMذD��)��?ۿ5�C��eP����K���Y���׈M��Gʖꡚ�<�{{��'f�[�X�T��_�z8quI!%��@�6g6�gw�z�`�~��%���`���ӽ���։�d�����#�>I�����Y����B�{�n�܀�+��:�з���=U�)9#��t1�,NO�r�5�v7�Y��ԇͥ��6�AN�1Q�1��
�e��qG����mW��� c��:-2�{uĬ8=Ǿ�h���/ՙ�#�dD�O���z:_0�2q0y�8��aT��.MW����<b��jW��:�=�*�+��V������ŏ� �j�E�l���=u�h�LL��l��rZI!i;������ɤ;��H���*�|����M�kK��C�߬G�|�0�	*گ)����b�-w*����<���1���h|ԻB�������102A/Q�}�� �ئJM"r����&%��9V��R� e�pl_�~xP�	P���ߴ���O��	&�)��N,�m?�7�*b4�Y�*wZ"k��c��L% (�w����K��º)v��u܀�Wjg�w��ٱ���R��J�	��L��'���6�ތ��^�y0	 St��͸�����y{��и��̇R�~BES{��z�w����=#x�fZ2H��&�����bV/{;�Av�I�����=K�Y)�����r:��2�H:��d@<��ŇjEԤ~��J�Z�Ѫ���P6�r\G�\��$Q��KXXm��)����τP�0�s{65��������������V
�`�	r\W�I���مw�Ο�4���?�VS�z�zU�\���x�gY��,�eU�m�Dݧ|�s@���(��oM�������i��ʰf@(-Df����V�� ���ч�RZO�3�c'
� ���q����O���]ƇJzPL1j��b����w+��g��Ik���>g@rM�c�0�g�`�'���ܴ�?��B_&w�����0�}r�)�M�.>��߀{m�&�7�;CVb��l�&5W_�6~\���
2�,d���fs��{Iµ�o֟E��u�rΜ2<��g�NG���R��癬8$���@�yb��V�E�\��UD���s�*���m.W���2݆�98F��)P�2�H�IÆ@��u����̢;� j�j`PC����^���SΟw�"����$�qp��՜��l_���OFj2��4F�>�[�˫m���I�	c�V3|w�X�*����DQ���Rf����������I�x 8V���w=Y�oM�:��(M���/OsH������
���u��MrUx��s�V�0!��^�9�S��;����5��-�^ [kr�*�xQ�A1;\ �W��ai�(C�����X�"G1<d��`�
��_b0��nQ8��.-� �w� �����%����U�z7.kյ���*&j�4=����};�S/�W��y��c�4��v���GQ���b�s�w�~g)��V���^gH�@nY�> $��d4�_V��]�NxW�C��1)�>�����و�y�W%����Y�Z]��?�f��$�&���&�J���:t��t\s���uh;� �S\��Qh읻N�lA��" �G	�"��֢V�6ט*��.g�S��R7x�5��Qa.cPfe��¨}����oő8Lk劈�a��0��1�vw�}�~2���0�_^�\M�`F�Lk�%�x��E���G�{��QY�*[�/`�mUy��!Ʌ��)~��e���ڱ�$CIH�.kq��\JF�z[l�c3�~vy�}�;9�I�zi��Ħ��w������RO�s�g��g.U�JɊ��=	��K�	@Ќ�g�u��jt-��"�}��3���S8�u���\��(As�>����q�A<��JeI�m�����bjK|O��uV�Q"���
��z������_R@@c#�L����qOĆ�~:�0-�:ֵ9�(���H]��:�[l�E^�^�-�*�?�#5:���v����1����l��o�!�ID���Ӂ�9_r��z}bB���� F�ALG�|���]5���P`K�08�9F�33Y��:�m瀙��t��X�:��#�\c�N���u�Q�:�çM��Gi�����(������\��d�}��gY���
;iu�F��^;R�?ɖs�߮�"�J�������&5G�'�[�N)�l���戤��y�ڱ.��Ƨ�-/��	��D��{�u��y����x(��2��&$�R�aI����|R�K|�d���ks^j�����/ ӷ����'b�y�h��^[�oSmS�s��Vq᠟>V���A�djס	
�jܨ��&'�1��|X�s�A��{�	��{ 7W��-�-PL��jQ�
=��=�,�t��apt�f55pTs�KUx�ҏ#���Ã�')��rȁJ��N��I���g��=�9�mmC��(�T�Y.R`�*�����,�z��ΐ)%W��	F�kD�����9dsZ_WΕ�?:B���F��t��LN�8�4Ϻn���T�=6�5���M��v����+���$��ѭ�+�\w?��2��:�4o�~��`l�P���F����c�a�s �W[�z$�g�t}����,�y�fӘ��_�5�3���`D
� (�d���s`>����X�u�����^'�Ĉ�b���d�EË�߈�]
v�J���1����>K���\Q�q�n֭Cj�ʢ��|�t��;���l��.�4�������~�@j����z�휣�y�P��i��tݚ;JTL-����3�����a�$?�9W`����||[A��d®�L�C���gh�rj �͇^��@8^m��s��}�~\�saqc6�K%e�lΉU�߹�L���l�YV��w\�щ[�Xs�#/	1���-��U���FN�)wh���J��ɢu�����*�s}e����T�J�[��O.�K<%��'׼��F�6�&����x��=v�S.r���&QՊE���6��9ڨ�$����A�m=/���h�;��?yRx^�x����vv��Mg	�h�!;^���W�_�'P�;q��5����#bG�=3��C��?4a����{�R�Ӻ-i�V�}Ir}ʢ�s��{�}=���h�8ɩ���ܩ��ZOM�ʯ�L7��&u�`Cqg�[M)��z_�Čp5^#�9޶ھ���x����l��w�plz�\���������0�O����O�ᶕn��k�� �eV��>g���ZQ�Z� �D��G�����v��b}�b{j�%��.��� X�;n=�h�9eח]ʢ����f�wh�G�o4��f����	�!������z)<����e��%�J���ϖK��Β�&�6ve�Jh�{�'���`��=CWh��jW��L�0��DM�xS���"{1<�
�3�%"y��i�=g�?�
i�C)W�Wމ��Ւd[�AZ�G����q����y!�	���f���{�N�~ [�To�#�`��3�ֺmcH�z3�p���^\Ӹ��0e%66�3G�珋x�ɼI�@���e�\��G�xt�sNh��'4/�u�NQj��Vg�k�NV=���6^�՛]�U��]�)��T��.�B&+�m�~b��A+���m�����e��"׬�0+��w'�N����������t�b���O��0'�y+4�݀^gGNt\�	� �z��}�{=��"m��#��J�qY��W��T`����U�aܺ�-��ի�덹&'߲�Y6Z@��2,�g�M�jߪ��	7d��c�2��[�1WIhH�D_�j�u	�I�=�{dдE��Z�p6Tr�Vb�ԙ���^�or�g39~n�#���*���aٶs\�1:��E��9�q��P�F�>�&׷):c��DY�����jg5��5{_����U׆�k���]�k�55���˱����]/8w�e�6�-�l��WcP�YW��%�{)�wK� "��0���@T�{z��B�啮������5(�F�����ĸb����ā	��uQ�[j��?�����Z�T������}��=���+/G�W�uk��e�.+��O;�	��k;֬<z�&a<�� Ed�dt�ӠEœ��A���oU�i	 �Kf]�X6^���^�����.���ᚑ�
';�;���=���%rҾ�r�{	�N\-�L~b��];���lZ���GM��E���O���#r��yyZ�O?#*(��([�T�=�ڸS?r�'|\����I��tdD���s1Ϻu2aBF��¥-�z}�S��UB��0LwF���̙�1Kzo�?��EkA���G��TwY���y�5ɖ)ʬ�]N��@��Tf���|"���=�e���0���Ȓ�Q�7��O����ǨM-/�����<i7n�?|[u��4�J�hF�o:jB��8�Tq����A[M���n^,���=����IR��Ubf��A;kʶ�{�g�>o�&��3e��4�v�љ7/
� Br�^ߺ����Y��}��yG���)Ϯ*����T~v?���˼����)!;�&r*߿*@2�/B��MX��'n��L���b��vU������%����x�w�^j���7�oz���7�V��:ߝ|d\��?���qO��[��\�4��y�n�}o5�3.����������ߝ|��	��oZ�=���d¾T�6u��I�ܫZb����p,�wml=a�\�4�ƶ�|���	亼�P��,cAK�B&�3rM�Ļ�HV��H
\Wd� ���f/A��D��4�	U�W/���]�^����d|�ދt��ٽ�ނ2V�h�6�vƏ�z����c\�v��>����萋��'Ir��T���ˤ(̈́}��9�"B$���~���P����u�}?%�6�p�I�� �X}��P���[�]N�o�e��ڃ�e�q�տ�C����̅�Iq�2-ٳ)�HE�<0+޶��p�ӎ��x�����r���a�V6����ض�k~ S�+W�s��J���2=b���;ל���7��>�
����ɩ߯~��v��d��#�C��{1���m\���7��TI#�5v�m��c^6��f�g��N�R�`|���7���:1T#�v�B��	't�>v������)�K����Η���g&���'R1�yV�o�,�h��3m�IK��V�����|��{3?4�uU*�ؚ�Ɏ�LW��&�����"�b��T��h�d�=f�T��E���{�qd`��C� ��s.�3w��a҃9��TD*��g$lSs�-�R��s���X�ihW�*A�dl��#���J��iW�J��H�|������+�N�h�����v��(@�Ɲ4�(�Ao�f�1��6�-5<AZzXX�,u5�%�o��;�B�قn�B�#v�����^���zۺ�<��&���fM���e���KsQ����dy�e��z�g�Ư�����+3ow$��m�ܚ6������ �<�'��٤��<��u|G��w7.0�X�z�-֛���F^2G�u[� )��E�>"�֯�t�k.^=�����P�B3*�-��	k�m.z?f�4iΥ���yǇA��)���-����zK���k�b�����obdxFC��$==�]��q�<<Ou��UO�_�7c��t��@W[���)H'W���2���Z��* ���%�{o(I� �6��Aݡ^�tѳ��uoUۇ���<H) HK7H7��twKww�
H�P�0t��Jw3t�tw�=>�������u�a�מ������k_���M�貦s2����_O�|1�h��0L	PO�I��G_l[X���M�jtV1���-,x�8@��d����ɷ����OTm^�0��.l�,�LW�����
K�����P�ݰR �����K�����C�>)�8�!h��u��Y&�kn�f�2�l�!2��Qg�Ha�#��Ȱ[��W��l,s\��3OhDٙ����DY��ww������+��B5���U�����%T1���~؆��OA�fE������*�T�$�1*{�벭�=7��������9q��
Ab�5�}���1�̒��5.���"ԅ?<���[�U,�<t�&�ж�Z{K�:-d}s��{�����S�`|��$���P;?ͨ���yz�ϱ�m\��_v[�po������t�/#��p��=���l9i�Ԁ8�1 (����.tF�9MU�����`2��io.+�R�p �)��?�SL�Ө�Vutm����9m+��1�sߝǍ����(E���d�q��^7c]�<<O������i��Dw|\�1&�idpV�F��[`��������}�����<�\��y�N|�F��=�� ԏ�9��H'_�9���#u�L�)�e���t�SdKV���ָ��K,�����;�����xEa�K��F��?b�_E[L�LF�5�)���U�շ쵧'ԁ�F��~�F�����j�7��$@��. Ay�|_I9��6���Y�.]9FM��a|U8��3v��l;����=�a&&��H!�>����B��D �A�P�1^��Z�Dm/�-&7�N�e�xP[��@��>GA���"ͨ4�2g�Ҩe�����9-�m�H1yMlt~����q�^X���~��*4=�^5��(:^��9Q� �0�XG>a�DŇ_=5��PGsځ_�YfVqv;��M����վ�#�����_�'c��5H4��1T8���UH�+��I$��3Pv�0�TR7�-��Dƫ+�q��Xl����Lu@@m�g8��Ѵ��bEj<Y�<E�<���wD��t�==y��:!�a׃E�z�(����j#�}�%�	���5O�3�M���&yI���Ұi�>��$�cF߮L�Kp�+�БD�`��O�-��>S�#����ي�����`e3�h?0�*�����,q�Ӎxj���l ��Vὃ �c�r���'0>�%����\�=���$��GX][X����K4�%��Z��\�Y`T����sد֊�?�&���;4W7��h��NǬ�V�{�ݤ�������������݄3 ��f ߗ�V"��XD�+�Ӈ�w`�yu�piӥ��u@e�wwb/Vܽ�<P�/��^}7���F��O��C��Y�imTwo�Or
�C�
�F ��;�x��TM�G�9���Q:Ę���_;�Ͼr��wB�.)��VS�'���ۏ�S�Y�/��s��"[���[�m�t
�������v�R�Y��+�0�i��'��G\����/2̷i�s�����f}�L��"��y���G�!�f��	P����w��/
G�����&3'�_t����3�����e`��kC����P�Og��ռi<�Ӛ�m���\�G���9��-�|Z�C���s�KU����&ǶOX�I^�'�m'O��=+��ՓN=y�t���`(w�+��
�>�ZZ'@���<��
;,W���t:M�J��vř��%�2�$��Ш$�_��z��D^�������r��j�G�?�_��jv���Qǰ��Yn�&����ݞ|�+�/ec��M#?+88p�{I�,����:D�Fba�i��_T�?�6�յ���̲�O��H@�*"��K�b݁�!z��?�W�)xF�BM��ݥ���� )*"LU<y"F�XL�����B��H4e:b4�$c����& '����˞ps�Q�lQ�䉂�Ϟ�.�_�����I	P������:��M���Ŷ癞溰Ԅ�Z��ڹ���xċ�.ծ��?Z4�/�0H<9?tüZV����7��7�h���$aqkR�/{2ܘi�_�â��I�G��H�Zy���
��s����'65��JVZe�H�l��$i��
�̀��RPͷ�ա�d�\g�LHg��zpM��z�VE��ߑo\Ȝ�$-uX���ƇMCQ/�T�֧,���ؠT�M�M�������Y[2Ke��f)G��*y��h�^ sN���C�*�W�((O_i�=��/����皹jH��M���ۏ�-|oÁZ�W�DY9��s�p�F i��hk�_k �XsG>(�V��2��H�1�f�;�4����8�2���i�Ԙ.լ�@e���W�RH�3�8����Ŝ���w*�Z� !�b����?��&	���gN�*o�zLΥ,�,�B�"kd�3�r��(�����=���vԸ�ׅ��4ت�E0*"�2*����T=* �����M���e;V��ٝk=S6��J��h3��P�N�T�E����H�H��F��d�]hx�JE�4�گt6]�AV�rN>Nh),Q��a��o��B���@��P�)n�
ӏ�.h���Ֆq&	��!PZ��E�C�LE�I�����&�N��HT�ʘ����@��k`Y�l�ޥ;�j��e_R�V`�;&�Pm�Z{�VKo�r���3ls�����3:��"�e�x5��V��/���:H#х4��� �Ѝ��̒�R�8�b����*b���$��"�Y*�̉Ն�.�Y�pI��Ί���9�A
���ʘ `X�2�<���<d�sob��і��1'�o̷��4g��=5C�Q7N�܈E����ʅ9���Z�(qP���P�Q���l4V��>�IOi�ZY��v+���Ҩ�`S(nw��bPW 7�<��w��vm�O�3��x�1� �=�!�LO��g���$�s�9�T��:��k��$�c��m�t�T /V+�M���$ϯ�r\��Ҹ�0�O�?+i���;a��}����
�C�����Ȑ������c�]��4��ԛ���:�j���q��j�0;5P`[q�T�����N:*|�?3�뮏N$G���8�c+ϟp|V��B�����X�t�㥬�<��N�cL��2l9Af��d>��plW�F\�C�|a�+|���C8}��>3���H���A��k�?{/��!U�(@���ǒ���6�궹��;��`��%F^A�T�Q*Gx���^Z~Z�9�e�3��$H�c��ƃ�x�{��uR]́&���9���y����0�Β�K�o(j�hl�@�g�f&8�5��2��6v��I&���7*P i�Y��TT�T6*7t��pа�Q��绌���<���273:����OP�4S��TIޱԕ�'2i-%^7����f�iy�d�]�4����
�=A�i�z[
�篟_�T��Ș\�gm�K���}J	�AAK^W{�64�9�Ӻ�[I&� QÑ�6�W�V�Y��/��I�gV����D��X��V`ƙ�ȋ���h}V%�8>��"iv��ג���`�eS�,�t9�3�)ۑ4��Q��3Vc����L�l����<mS-Dꛦ�%>6p��tܞ5;��bf%1ZFX:�.ޚ�s4k6��}3�6�7#$9hqVhЙ��2����]�+�O}��(:t}�z5W�}X��~��O�P��,jmBV��}O�mWr@Euj�OwD�u��(����F��m�)��KA����$�;Z7�;��>O|���@�	����̾���G�tO�`�����'E� igZ��*����Co�k*�����2�_�l�i>�}��w����o-*��������\iY-�H�n@��끥Cą����M�h�7�s��I�$�%|�/������&� Hb���Q{�J�vz��?i��cS����D@@m.��>���wI�����nN�S���|BE�����Z����0z�>�+�i��ܠ͈�"U��GJ�Z���5���ߛ���2��g�\����G��]�	nDt�\D"B�ˑ�@�H�%S�׍X3��� A_L��3~[.�(�+E�-��!Y�$����v�ć�_�X��~R1j���a��\/W�|��z��TUd����I��V�G�	#�	�(M.@Գ�g�o�4ެ�c���-�d�e[���2�����fd&�>"e�b��hz ���!l���H9�K5���4]?��3p_�5~����Rm
�G�o���pkl�0q&?<� 1��|*��\�HAE8Ŝ׈M��#��C�~����)M���z��Z�d����Yv^|��s�T�{���RfgDqJ�A&�,p�_x��8[���}�˭Kb9��%�d:/h�MXG�����)�e�i��e0���T̮���Ӳ9���Q�2��y6��ޘ
bT'���Vnype�hA�,Rk�߉�L�d!��H��sq8�d�"FZy�Aa�E
&;�#t~�ɗX������4B����ЦC�}��r��U��x¤�,-���D��/G	u�jW�|2�����^�ɤ�(�3f,Os@�o���S��4\M4j�p������Y,R�,ET�pٝ��i�i��w9>C���%���b2�U�N�ss�hj�k�
d���v�PFN�#�:m�z,Vnޮ�Q�@c���<9���+Š-Pc=�� �Ԓ��
���-x2�^��i�A~����WF� �82j�F@��5nr}�W?��2�]�"�{����F�hܲ@�����m?w�KBۤ�~�8�����2�!�+��?�g����
��_��"|��%rV@�7Kڤ��>�~����S��5�C�(�~���s'~�cÊ$���F�!D
�'��y�ꮘ��+�<�6���������޷����G'ֆ�7W��ɿTX���T�yƊ�2�5������N�� �C����Á΍'�á�W�?���������A濠:�o�b��L�ģ�zU�����1hb�*�_)��v�(���A��ȕ{�ֺ�`���"�k����`/�j#����bOQ�ɚFleJ�Εi}U��M����r
	*W��T�	���o/%o�w%"�'����\]��ΝOn��a'Z�X������r��[�~��Kp��ȏЄA���'�XK�iɡ^�u�E�|]ӛV�"|��n]�L�%6�㽩�2�9���N����4Y�T�H�|���AF��KYx]���uc�����C׽�����x}U�)�Oq���'K�&�k3 '~2ޥ�,w���ߙ����hUz��ף����x	5;��uہ`͛����5r��B��՟B��ŗ+"y��O�G�>~#D"���{�%��CP��6G����#pW��	���-벏c}��M�k�>�{!�H���|-���-l)+���ƠT�v��|�8'G�p��:����`�UN	lwl��#*(�x�Þtc�M���2ތ f����>�z:l�.KY�	��x_�g�͸��m�6��u@��U�����Ȳh歿�5{���=����py�(]ŗ���4�#�u�q���Xc�D-*�q��q�}$�n�4J,/ݶ��B4��C����v��R�W��3����S�^�<'�;�3X2�+p���oket�yH��rn��j�N���8�L�^���Ѯ��	m�$�Gޜ�p�mc��A�+/:���O�U�o61��,jv���l7�=dZh�<�Ke�J��M��)�A��V]mnr����>���O�|k&����'7kF�+�6^����A\��.��e9�ڒ��W���r�4P�����˵_�߇�Y!,�<���\��&X�SK��޴N1j�d�Jr\Bp�I��*B��<+a�ۙ�|D�i��z�^wfQu���_�p�3���-�7�۲��c��7�ﲌ���F7��V��
{��K��
�ۊul���MA��\�KA���RYg���	��|��֠>O��bNR�⾐M��1�U��l�H��x��20ͣd[�{\�k�;6P�F��(�0�?Sᛸe9��Q@��Zj�-�ל�zD7B����T�l��8.��,��0�^?x���P�M�^,o�$����T���\o�#Sa^/������n�8�/����a��S�N��x_Sk5x�mju�l�8��OH�$ϷT��>�|��.�8��}�4��z4Tts�_[�~=�8w����h�(�@��;��
j�{TL�]�s@��ҹ�!np[�Y��r9�P3��japor",c?���l��VdQ�W'�}]�Up����_D�Y{�){���4��K�?���[G&�m�Q��Ei�=�.������C�����U��8�H�T��:?ŵ�}�	�h��n�>d��O�Y��y�g,I�Y�}��4��S�ƄcC�9��"��ZG"�Fs�^M�C[��9_8��{e�2 no�P?�Xj7ad��7��e��Bwz��c�L��0b4Af o����6r�5��s�������װbR[{Vx=b r��wx�U��ר��SW�1�:���r�58�9� �x��]BNB��u�O�O�4ή�\m-T�y0T���1P���b�vt�������Ή7��I3X���k�кa	X)�	TAW٥���u4A{+M2�_�>�շA@�cz�p�2����B>9�>n��^�����e:�J��Y�3�of��4.Vo�Mp���Y���64Гf�eN^�,�<_���0Z�۲pٲ�M<�ڳ(R�`���~��!�X�ø7K!T�Ӛ6ɜ�
h���Ė�|��Ä�l����t!@ߜ9�*�P�xl^�*:�*�e�����%��uZj1���esw"i>�ua�@��/I���<0o��'�%D,��.VF�}(�~�Ί�
�~��g�^�q��x��r��w��C9�!EWe>���|�+s��YH�t�V� ��~�1��	�iόr�\��LF�%J����d�p�z�OUJ����Y�k�=�F3�m�+���)�sPR���M�����	Ķ���%\��%��m�/���3'�N]�ނ:�E\�a�Jg�s2`qXg蠫C�/1օ�	�_�Q�r@ҷ���N�Y6�֯R=�a���L{��l��[gY�=���E����?�͍(�/Hh����' k=�Z��υ�R�T��>-������	EA4��}��Ow��(�������y4�@~&���z�n;�������5%��1{J�$���z��z��Ɇ��aPMO�:Z#��y0c�ʨ}-��O����g?��C�V�ʒO	4��g�rW��� p�`��V-ߝ��/K�������='f�Y�*CM��.��t.�i�v���\[U�����p��as"bXGꦃ���N��4-�����0���6���5��aПc-���������kh�����/_�G>�p�����O�bƜ�͙��>%Y�@��{�k�.m�29���r?e�Nw!�<Wg���"�����X�ϒ�����C��Kz��S�h�a�r��ak��� �&AwN�ڔF�YYX3��y ���I�p�U�
�Nι��%'G�?g�%��D3�u������L�O�It15��DiN�H�_p,��X���eJ<��y�����B?<�:���mc.�z�*�e�L�K��W6%m�Y:��_�TX���O��Ͱ�7���Ju�0�@�d�JYV�3N(&���5�t#�����c*N�K+��s��ZgS�_m�&Q�AH�݆	c�'o��ﾳeI��;n��ۧ�}XO�8�@~%�ױ��|CB�*Ո����LfH�Qc�#��[�E���T�?H蓬\"b��3sww?�p�sL}ldG������L�ͭ���R�����#6�ĵ�Q�!�:�V���0W3s�/��d�w&0���נL�+�c��!$V&{��;��`?�?-?6T��6�rh�p hU�A�CW>�j%ޣ_�ᅫs ��G^���z��l�F�z�QH�>�9y���X�8B�WmI��{�����Ta 9�:�q��|`:/Wi��xF�y��۹�@;�Jݗ����a�_"?�3v���UM} �4��4��	r��ɪ�'+���J5���[�(��G1�d����َn�=C�nb���K~_WW��TZ���[,�@s������G@SI�gS�[]EԽ3f��{.CG�ڹ�FO����0�;� �q�����(=����:p��ll���9%Zg��/{$D�� �F`��cҀV��u�D���<����to�yk��_�a��@��l�&<LFK"����B��X-�u���9���L��}��)�]~���w ��;TXϼ��v���A�|���漸�p�%��Xa�ao�@&δN����e
�G���8����<o�Q�1�װ��F����&����2r�ȉ?�����S����_�h��A澰�Yt6���=����p�c�ᖪf��
ew���"pJ�R ~a8y��
���\g���4c�6�$�
��=��J䚰Ws�m�mt	�G����u]=6=)�M!Ͳe�������GYAf���5�ԥ��.��RUѵ7G�
�N|V�i�n�Hԑ�uW���2q
�eC;3�r� 턃���v4N����=��܄��d�Ĕ�A�AUU:����3
;��}ڼ�y�Us��$'�N�4�Ή�{q-[W��IGњ���F�>�,68�fkl��ل����l���W՗j3~�q�9֖;�����k�6�0�F����__HU�]Dw�?������`�:�_w���B��3Ieѹ�@������AQM�Q���/��G��_��w9����'�
ye���ŗ�G@5�*5�d
*�}

T6
���xI-<� ���<��a��e�������:��k��ٵY�]hH�+��(n*ֹˤ���� �?��[��)LH�S��-��&ơ52�;�(��I#�F�q4�t�A�2�Ib9���ZU"N�$t��W^����!G�$7O.��ڛ����E��F��S-8]��3*�	q�C��X+�R��Z�rY�E0���p�L�JMGQU�M�,��L�}T��ʁ=�b�fO9+g�Z���l�����(�
&�<��O�=�߳ ��%G`�Ԙ�Xj�o�ܴ������!������4V�#'� ��ݓ�^�7�ޗc�y͌�����r��KN��Qg)Y���y���ɲk�̩1�x���x��cIP��Ub�d6�����z�F�ʆh.��ќ��&Z��s"&�ӄ�0o��V�ǜOo(r�����ޮ���hX~�>S�D-laĨ��<��Rc�G'��s2;$zۏ��&�DF;>�	�:��f"��+�`jV�m<�-�4wQ�^�+�,�D8�i
�Q&s �b������Y�#'��si�2���TvQ�?~e���S9�u�2�`�������
�$x��S�һ�5U�(ƀP;= N��2�����\�T��o4�Si�5����������"s6Yf����k���J��
Ҫ�v�iy�4���Jn��s�l�HG��\@�]��Ո϶��f�D
?�����!�Y6_����!W���׊����S-�'�����������)��2�ے Q� �Z��|��Qx�
�<k�����0��q�ǿH����*Ď&�rn�Q7@uT��O-�W��˝������@Gx3y�!=�i0���58�`���u��?���+�]5�U�k��������+4���ݹ� �Q���8oSS�m�\���Bؗ��8��
�%��(��,������%����T�hx�J�0E�D�Ϊ�KMB��..�*l���.fq�煓��8����_mf�莚��Mb���?�``8�����g� �4\��|��䓜I<�vCc(r��Xu�Q�
-�'z.�S�KH�6}���C��[nw~C�'0���#�9��G+��P�����",�bF/`nR���~��|r�i|�vb5��4�ܯm��G����I��SHfi/��g���/<���
袒<������G�F�ָSkk7Pc�|�uW� VN��<���)�L>/Y5Y�M14��J������ύXˋk͹Gӥ�@��7���Ao]������?��s����p@��G�4f�õ�݂�'�ͧe��Ӝo=���ΐ��!�Q��F��߰L���_8��~��>�P�2l�RՁ��jK�Ji�6����A�[��h�*�w�s��TT������ͷz�Y��q�*���&\����&4A��H�i�^��x��ܚ��1RͶvc'j<9�D��� �zGˊd�[����,M�+o�J����6�=e�y}"WS'T�J�&(�I�1(�")Ws뇳�̧Ó�,[\�����(n���ZY��u����\M�6/N��dM<��X��5�˔w��|��f�jNV=�q�!26�Wi�Z7��c�5�n��U3���8��A�`�Kkcv���O��JU�T�,�9��������ƛR�Q���*�n�FVj�s���L-��d
���.cR�v$8\�#o�ih�	M&O3G$Q�XYڹb�ş)���Z�S�pBh�z~m$&aN"���x�Osy� {�?����x�J�+�hO������o���+�)y�o��o�ׂA�{s=��K	_(:�M��\Rη�m���O+�cF��y0�`d-sk�a�r��R�vu���B2d��a��m}��N��X)2Y_ �WstS�����|�ϩ��6�/Z{*�:�X�e�Qy[Z�(j����'��V�N�o# i�q�'��O���^���֮s��pO�8�Vr�LYI�$�[���͊Ӥ�{Ӓ��n�*�~[��8��hi�!/��>�I|{z���.��g}��!�8�q�$�>=�g^���f4��~����^�P)u�bKT@g���P�X��C�y[}���L39�ss" ��H��DB�m���$�{��g�K�\��4��:<���tW/C^��\��V��fNa�K��\�zz�@�<.M�l�z�nI6�8�V�V�$O�D�Y�D�3;�v�*8���^)�=���瞱��30�SK��Z�i=Yp���wc�Q}kdn�6�<ƶP�r����C���g�m�������ށ� g&��޼��1�	*Ei�ڳ�,�CR���M���O�u1��4Dm�z�Dֻ�J�ȮG`�E|��,$	J����I���#>
B�Ӽ>��6�%�"��X���L�/�(�fj�3Y���G�rȝ���=��H���^�����0��WPƀ�TGC����a�-'�U��I�~�6|&=P��<2�JO���k�*Sl-�oYo�:�1-���g�Ë��o�q,�sR��q�/:eK5��/�8:fT����];�9#� [Z��K���~�#'gg��ƚ�>gM�dG���*�C�*�]������Za��a�̐��{���_GC��W*�����:�<�%�u]]y���;v�¨�|sx�UvJn�B�1WH�3��B.�)1��|�iw�mZecYٰkN��
�O�g����Yg
/م�>F��_�B���:����]�Q	�f$���[�X��F�,���JY�":.��R�Hׂ;R7�ńL5�����QXi>P��T�ԥ���j;�,B�~�����g2%���b�1۽�w�m����#y<O�J�l��L�|�xBz .$��~� ���/#�x(�S�ҠS�=ӡ԰�W�}_�Ň�[���_���?�R��Js�,|^��_N7Ê���B1�vh�P�1�xQ-��c��Lj{{�T7�"�� ����B��;/Dx-'"={ڬ�5~�����5�a�:�y���|�RU����1-P��^
���ZYzn�as���l-W_��x��t�2�D���i� ��H�0I����P-UF���=	eS�.^d0��{�������֯~�y��BI�
��"F�R�C�����^�c=�a[A�m��̕yH�g�ÓB(�,? d����4��}�#qGi|�~5�E(��6Cw"��D���%6��s��Kx��N�<�{ӈ��'�2�đi�)e����?`Mg��o���}S��I�-R��_'�K��^��y��=r*�J��e}Эv+>����B���z��Ja`y�@4�F�iu�����2+,�����S'?I�wXѸ�S��;�r],f;��"X���K�L��<��ʲ�T򹾥m�V�z ��u��|{�,�W���a3bF����
����C���sxg���W�=2�I�y�P�t��wmd]*�`>�QビN��.2#ϻ��w���-4�;�w�@�>��Rh�n�7�Ƌ:nܼ�D��o
���ڌ��m#_�!WW�bI�;ޜ��MX�6VV��'���I�������*��#�4�$K��-�� B~�b����H����}�(X�WmN$z��6�~|t�c}m��a0~C�ƶ�d����'��h�g�#QV~���Ă�x����5�d���>��L1�jkG���������仒@J؏,��� K��̓ ��\4P�&�S��[���C�_y����~����G�������k�Yj�N��vR�7���;��c��*�ՙ_i�ZoY)GD�`C�b�|��<�A���"0c�[�GY W�������h)�=V'(8��nդ��B�?U��c�ݚ|���[����������:�J�v���|Bo0�b2����tS/+�u�\���L:�q�g��^���R<��.�T��]Mb�Df��;�Z%Dl����+!H���)�^c�Fۆm}�G�����xY�V�0��҄�XX5��$�t�y}�1�R�'��i�����	������+�Ƚ���MM%Ѳ�(^�($뫣L�̍׊.p�'�I��41�����2 ���3*��'CS
����>nE���(q���G������Q�%�&}���߼)^&�q��x�J>ed�8+�vm�Y��j�U���	�YZ$էJT�$LY��y{n`�6M�_#�L����>�SK���.]/��O�bTp�|k�G�N�}K�Q���p�H^�eġO�����ָ�?�a���a&���=f�ۜ�:�u���f�ïg�*%���'}��*��|")xN,M�y��@�n�T��b�Oe�h6L�����F?�KO���w�
.��?4V�`�RU��V� Rȃ쪞��?�JXx��P��4��s���'f��7�x�r�Wq1-e�
�p����56�ta�y��C̝�M���L�c.�6�M?%Hk�!�c(�A�2����{i�z��2.O絉G�c#T���f��	��	��Ji8��a����R��c��# $�3��X!���'���_ض+���S�%�fg�g:}7�^��)b���2�_1�ĕ ^p|��cƏ�/Ky��S�d�t2GzX)�Q�ۏ9g7;t���S�SR����@�&Y���3�ː
���	O�녴�064rv�c�X����P��|;P�uhi���F��D:��Y��,�������j�g��&�LVyu <�_j�KA�M5+�*��W���W�j�����I��/6������=��KzH��FKK)� CK���/�+zi�:�@��qa��f�ѕ���6��-�=�F���i��!)H���S�$��>����E��)?T%_(q2�er�29ry�J��L �D@~�2�G�o($X���|�WB��/B����ށ��͒�Q��^Uk�(�`F%|-���&�z�}Ă���Bk!��������NTdMvt�p�>}fً�s�_#�)�������9���������I�����*@�H�z�R�"�5���C�F;�����68+p=iډY�#L�dc%�K������T���y����w�p��MzP�t�U�+�)ӕZ�Ck:>����~�k$�S&`s�ZW�g8������Wv�	�o��3�b\)����[��S5#��2��]��7@�дYD�yn:�>�(
KI�[�ٓ6���88_-����%��[qE��`�N>W%��� ���'ҾhX�)�g� AOۏ/P��>��|Z������%_rk[�^�MCS%��H3;0��T��=�V���Cf��v��e�������߂ä0��C@7�aD\��~QmM����-1˔�WY��I�,犢�����Ɓ������oǚrx`��bϫ�7<�<�*�9�w(�`4ྷ��0<�����"�?'�f�N�2�ܟ�Gm�V��?q�t�ò�JO~~*N)Q�����j����W�k�w�@�Bag�X��àF�o�F8�+��n �|�5I�@�X�e*���_}`<�x��|��
 �����f�%�?�ac�
���|8��{�)��րV ��
ߟm.�{�mg�����E3��E1�����;�(��n���b��T��bG��(�/z�������t����E��n_��OD�U�*r~q7��=��v����<�B	6�y%z��L��[JOn*"'�~E
2v>jL���-�?1���`.����0���o��7�8�s9�^��,F��IR���DA�W�$��0���G�II!'�7��&�������`���	n�:��d�m�U�R`�#�U_|_c1���1���~�� �7�4CψSBѳ.-��cc<�Z�Td�JtpNjBպy#v|q�.��O�����ܮ�
I�(��G�U�b[w�&�κ}��S*�MZVAQ*��*�6}E��3� +�ߜ	o>���Q��[��ֆ�I�!#�Q� Y(�8�G$���7��i潔t����r��A�R�oj,<�a�~&�f'%d�B��A�X�,�9����t�9#����z��z6Jpڔ^u�R��aDx5OR�'�*�.!�;�@h�*8Ɗ.�鐤43�a9ƟV�,�
4H��N�Rm9ݎB5R���~�qA@������خ�Yy�����W2ڔ�B,c*K�$⵸�-�h	��:�N��
b�MިA>:8G[�����BN������N"R'`����]��ӱ��&��>}fF��PL�����M4%��&%,Si�?T�H\��в�\�]�Q����c��Pʌ�6b���0b�v�+��P�$JT�v�Hv���Hm�)�K?��e ���Kl�ٙm$`�kKՂ���߬J�)φ�G���\��.�2Լ D>{S�2��qze��!��Z`��"_ y���y��|'Z���]�	�ǉw�BRo��+�ؠ���Qe1�o�x��`�#��g�t_R��̦8i�5���D�?��w��]<E�%�m�uT`���Jk������T��;c��d��ۍ�a(�M���&�;�Z�bqU�`	�$�?����?��F2]�~�8�t\��ڟ~�R���i��|N˴]@p/Ͷ}ׂ�4,��K�����i��� H��MA(.#]~�q���eS���	�Y�G����ͱ���m�z��"�qҾ�<�) b��ڃv�u'q(n7,ϟ�~-͏)*�KDX��e��ntF�X@	����쳎ZPf/]R���O���&�DK��õ�h��<�'\��#g+m
�<s�f�@x�e�TY�\N�Ӵ@�߲D���Q�"�z��O
�sڟ�I�R����z���S��k:0~�JD�uDL?jg�Ls:�%k�$� ��.J[Su_���}�m]{�:��e�[�;�T�������D�UIu�4c7�H�ƪ$��|g@w�� �t�rE(>^���v[�E��3�PH��>�������V~��ni�hNݪ����y;Wby��Sr��1;��g�|!�3=�c�V9���`�u0��p}�')~�Xw%�1B%ۨ�zOw�<CɊ�b�E��rG7�"Z�dt��G��'���\(ET���}��Xh��v
Z�����gi�o�Q���cדh0�xE�:|����L�,yH�ŭR�ol����x&<v$�SF}�Z�ܮ�BAZvwWnQcj};|���6S(Qs�)V�rԷ�!��`�*�4K�Z7WtUy�Š5,�fm�/W���G.ǉ
�
�nϡ�%�/��7��Cc�y0�� �9B�J/�����&�d)�8=�{�`���~*N�����x��z�{�E�Z!K]�p��tW�%�@a�?aKX߄�_e��k�?L]6�
&��-�	9`������	ߥSq}�b��s�e����j+;ʄI�W��M��%8�ǭD`����铨�p������5[�����
C@3I�8HFn���u-E��ֽ[̓�}�6V�hGI���d�Z�=0��씞�Q:����y��*���"M���)8��w�����Q�i~���f+&�5ᔞ�M:�޶B�\)[�ap��E斛Um�=>M=�n�`�uӰ�R	�Lw�E��>j��2�]�~-�c6P~����\�0�ޝs-~������EQ�'���.��aWpR�<���U2y R�'����=Fm٧���[�-A��oL&����>�����l/r�[~����Ňu�n}���@`5�r��t
ڈNoj�V~�����<Ox����'���K�;xap�K��x�U��6�?���&mB%����&3��\�Kg�'|{�C�P��ߣ�����2�tj���6z7+1�s���)�ĭ�i��&�1 �,���:qXM���ɼ,W�}�w)���ȴT�Ō�<�х��#_p��<�����C
���� 
��y}�j(Ӳ��G�.�?2�y�{�2�X�Z��2̪�P	��\�0n�"�|e�,�q�IJ����?w�� eY(L��.��$��ǽ)���H�AJ	���*.fx����OL�g���	m�c��]�IL�o�
}�<�b�4�^\�s>I���l���s��2�=�Y4U췳��ZEg�'3��|��m�E5�a=��I}}2&ڦ�5�)�X_)�F�y�VR#�j��-��ͩ��N4�vR�7Z�_#V�K��d� �χP�j��_2�bC�/���yyyC�.��\�!&t�*O��
o.���1��������Q����pw�q�x{�+�g�]�᳀�7=�R�S�>�jK�7��ƷA7x���f/��~��,�ۜ���Fqfh��|�{	�Q��%tg���I�%��HI2l�~n��5E0���� �L���j�x3v4ut�1�E���C���q����Zn��^��q���Wz_�6�<qeҒ��y��x���	�.�|<�	��.�c����ۅ�h�P����U�׫���M�����R��R�:�0ٮ�H m�	wλ�f������Q�;s���{E��#Z\���RW��4{���2*���@�W@�TA��D���R�A:@j��k�n����CZb��{f������vם����O���9OG��Mp���Ȉ��.��C|V�C�@�+]��2�O�@4/�T.�%ʓ��#��{��#��Ie[}�����t+>ޜ{иD��m�p3B�ǧJh��������}i�����Hltk+2Icw���JT)w��ܙ���'����-�M僳)���O���\�R�s���ύE���^�;׭P|�'G���:@���:!���gZ�bB˒[H����l�t�%~#��oep'��d����j#��m��M{֔?7�g�gz����[��rc�m�����r����CL7����� c
�k'��
��ٛ��+�'�e��ʯ��|�z	�՗��H"9�.�
E^�k��$��_�;n��tre܁���o�eE����[�BK�rGo�o|��w�t]�B��(ݮ�$|��׵�+�O=�sR��]r����]���ԿKW>~Nn�������=���.��٩����lGH���H7oR�����o$�<�_r�t�B��iBҨqS����bC��';�rZ���e�R����W�7��c"s����}c �.�1{~	�yN0q�[:�7�]I�x���W�����FW��+�M#
�����<k܏�8��utg���G5f^���TF�c�.�ď��Z334���/Jov���V�vQFT��f'��Gn�Ӆ�mg�J�w�l�dmy��\����z4��}��2�k?���XY�=�c_i�+�ڱY���}m����|]g/�՞;�� ���&��u�\�d7�|�MKQB J�k���#���'������Go9�q�|to���ĕ�cD�a�`���w�"?O����8���PO�A_H!f�qP\$F�Cj����s����^��!ڴVS�]�h��L� �����Y�T���bc���3�W�͹�+n31q�K�;����i���"��{�,Kbd��
�f��v��E�����s��R�]���S�y�����PX�R�%���lMc�e��[SNdg84��&{�(}/݈�}}18/4s<��j*�cS&^7��A�	��pC� q����������6ax�}O�}�_ꇊ���Ϣ��d˒��������+`�IH�G`��[��r�	ӫX/j�=п8 ��ˣC7�s��?�������ţdf��7��_g6Г���Z8Ӽz<B�~D��6���\�*�61[�������osD����� �h��:���Qs	�5�j�+��J���sb�z_V5�>"g�l�#şz��F(�P���)q��#�<C�H�6���A~]���J�+ͬ�}��cЃ�y]O�ӂZ�!��Lwǜ��/�݃߹E��4��'Nʃ�~���@��S}��4���}��rl���i�`�尺yv���{��S�������I�O]�#^�]%�f	�0�l[nR�OF~X��.��e��y��/���g��8/"&�˒�뫠�����f�"����6l��,0Ύ	O�2z�w�Fxз���f���Ug��׮~��̎
�� ������'�mL��)�WP���ɹ�]��S/_V�i�s���Îٗ-b R�^"$yrF�1�{B6�:���w�L3� nn[''�1����ˀ��аگO�Vd^6��F(��7���H�9�� �y�c��h�^C������������ÍZX��0KZ��?3��5��u��IY>�x�!=��
�0�2�l{�cu��=G	�9ߛ�D��~*�4���0q<�??ԧ�j@����� �A�/e �'v��~���#La�P�N���݀���x��T~���0t����5z����/w=��qy���5�z��"�6~@�L�Mg�4�o�^qM"�x@�>�����g������#��Z?����?�`K��ΨLS��X\c��*Z�&�tl {/��]��
����j��q�����.�[�p�hV\��ψG/�A7�k�nb�銌Z\>�t��6�N�¶�^8��+�轢NT�������nS����YKqi�"��:�6�Tf�a�4֫f �ׁ�O��h����o�\� ĕ/�:��쿛��{�I���.�?�y#u���5���w5�tѷ�GJgΧ�4��]�����lu�;׿w���y���n٨E��!�?���V݊2޼�v��Nr@N%䛢�lD3����L�%�F��:��#���.ˀ6N��D�p�BdX��6�7��	�q�0�oj��޽m���w5u @�kt��t��[t'�+�.���X�=��Z�.m�ȴ�k 	�w̩�@a��n�"����nJ�t��tJ=�[4���*�Y��<��> �_���gN�`�.�i�m�@i;��|y�����H��]y�o�O�1��qy�%�r���Y���y!F	;�
9E�|��������Z~���`�o����y
�Lە���[ټ~D����J��	�C���^��On��ɢ�eN��=����ܣ~��������[M��"/�!�	��5�΂i�k0v=�FB���G
����Z����m�����p�U`9Y�?����g�%^���Mu�&��n/ʘmG��I���0*�| ���z�����d���pM��`�@�(�F������ƥ[�౟J���ܡ2B?��3W�5�I�ern�i�� ��2�ٰ��tt�>�Y�?QK}��(z��VwNl��J�G@���dC������|;�2Dv
�)&��Bvd3*L�,��d�_�s@mNx�V��?x�� �=��ۍ�l�';�����9�����A8��i��o�ET�@M�����ő5��̣�mB7�}��]�ݿ�/�8 �cع><�JԚ�@����"�c8�2-O��OZ0i������)��ikb�ʬ�-���2-_VC�����j�*�D�������V�M��V*��-�/f�9h���$��j��
G'jϾ�g&�Zeƺ
h0ꄘ��S��c'�.;�Y��ؑ��T���n`�.�"r}H�o�RTƁ��++Z�}�I:5^(�b��i��~����B��`����Ǻ��ɘ�4�ȶ"�B<�d�Y�0��G�g�Z�����E�mC�4�-o�'ui$�zZ��!Sf�������i�m�S#��v#��kg����W��"o�]����l��;N��+�W�x���F��'�f$%�� a�$�_�/)�8�3�4w4�[Ȅ�T�}��H��ѱ�F��{4l��-ג���Z�A��̯��62��Tߪ ze ��N��0�q]	y��/�E�C"䃎�рO^��V%��D&�A)���+��!�R��u��2�_�2�Je11z�h¨�K��}dT��}?$c���+y��!c�I��!c(]e7�I�F��ȍl��lm�Ѳ5ߊ�=S���B(���p�N��W� 
@o�a��	��� �E�$~Q�v=umIH�0�?���q�%��������[W���b��#	+�]ܭ#UOF[!��P(y]�7��6�lR:�|{&�O�`�E�ĕ]�T?�mݦ?gI{c�f��`X��&w��$[x��= �-2��^TQ��s�&ɀ�����.�/#��|����$\~/J Ք3'�+��>d�`��y�U�-64��Յʿn��_�M��z������Z$���H�������2)�M���������rBO-���d��I�����~=t��P�e��~�6ӽ�����;�j@�d��?�6q�b����M�^���`�!m�]�Vy_"4I'1�,�靹�⌭�F�8[�]����#|e ��,��)5hb��ݬ�g:+�T��OqЖ�񃬋��KG�7�l�{��;ڳ*xq�KP �7��:��Ђ
E��<~�/2�'D�J&�n�w~ ��ј;Y��Ȳ��Y&�;Y������ Y�]��l#&$¤�f��f��9���h ��U�l��!�?���(��hTxT����ia�t�� �$n����:����y����̵�����M�usH�j�H�!y���.b���jܔ@T��A"�@���Yx�}�٪�/BD����9Yp�@��y��<xH��Ș>zud,������Ї�_eE�/�e��9�����wi�u٭�?9���ʞ������-^<|tִ?Lm-���n� Yd7�m還�<��
�KV��>R_�p��E7O{/q���Lu;��]�9�c/8=S7��d�igg���i̼���X~l]Y����J�'������T��W��^'7�7��̼��f�=ZwuI��ƍ9jbp�4�$�r�YZX0��HO�#���� �+���Ka���lqײ.o3Ύk5�� �҆��-Wj���rG�M��KP�a�ҝ��f#�YU��\�z�CGٸu�vW~LAfY�F�  ����E^��h�f��ioJm��y��j8}x��ف,�D��~��;�x����齹�W�ʄ3����@,��$�6�!�/;����Zg db����O�a��O�� N=��]����V�������r�3�ٿ�����(XW\�P+bG/Y1��am}f��Hk&�3}az_��
TUT����n1:�ߟ�TV<��a�jܸA�jۺ�=���ļ�(/n����[w�L��\��n]/6J,f-V�� �9�=������kZ3����e/�"L˚��"�6+V`z�������G�����UDG�%���?@L?8�Br�)S�B6�>J�o�>����ѓ���CgȰ�`V��b?�o}�c��-[xp2��K1�g;1U/�?6��� ɮ��|k,�2w�!ֶ�+���aR8Lp�n��^�t��h�c97��J��9t��w� ؕ��������x`��\0,�|��)��I#����l�]eR
�U���P��l��%y�`�̮���+�M���M�g2rҶ3z@[
˪>�9�����v�:m����H�l��P��Sڔw��ji�5<������8��ݍ�个ڈ�;��-*T�3p	��;V
�1kE��Ykv��m�Jx��m�Ƞ,=ۈ��_艌���^Ԭi�}����jDA��~��U�a��u�tI����pȫ�ή,)0f������D%`��pXZp3=oxת6�0��b�O��e�'^���DvZ$s��:2#�}TVU5���MR�џ�x��z2O��y���{xw��E&Q�;�����e(+�4��]�3����6k_ǣ+��D;:�U�3H�L��;���ƈЄ?��e�зOx�W��_V���#Tˉ��<��/�ʫ�xB���L&[��yx�^כ߽Ʊ��L����K4�n�&'E�{Vbm `�8����ʒk֤5'�{�b���f?.=6R�ݷN������k�mMd�s�S�˙��6�r��9�1+y��>�S��s�׾��,��>l��<I	[����YL��ٜ��}G�<�D42�
�CE�	t��2��2�����N��z�4z���an7��^��֘�Ƭ1����m+�EI�:G[�(Q�}�
�Q�*X�M$*�Uӥ/���\���W��]��	���[�5���?5�0�峏%�IL�����c��,��&!�tUAHPb3��nD����.��q"s� �>��*��|���nK�n�����x���@3�쬐�a�%#7��f<�����5���&�]���c<��D�_b/T�p_~`7E���@������ѓS���7ݍ�؄�)Z��j�:_�%p��v;{l2�����ٷ�
fL]_w_W�А��x��Qq7U�f��N�9�ti�P�5�]��%S��O@-5�i	um`.��B,�%�����24]ƕ����]��F�k:�W����v�C>xA�תm����V������P�9�������������K˅�Y�����R��{�x'8&��>�&[�%ԠxF�Jl�	�Y�BdL��aEE��Ƃc���hw�L'��8�_�;�G��e4��%�^�M6D�R��'Y1<�*3�H{�ͦC����6M\����Y��D�R�nZP;57��M�{�a���^R+��u=H����D7y�,���<.�o�����40�w��/̼usLS �L���4p��`�E[��x�=�-�F~�o��q��4���gx	�����c�"�bH���[ͤĨiA�wo��'Q�o#����P#obJܬ�3���L��|��<xӗ�଑U��K���e�&�nn�2'۟�����$�.��k�Z�Cw'��TΩh�Ґ�+a_�r�sq!o]w�9O����squ��$ֶL���y���$C��TS�GQ�D�PO�:���K��t�֦��}�Қ�����i�[���Y�h�Yڠ������+������}i-��P��sG��}�e�5S*��E�G���H��z��JVшfބ���Ǯ+���r�����#��>��AŞԝ�n?��trr���n�V|?�A�G�x6lFЪ�Y	[ޒ��CF�MלOפ���S�4g��D�fS�b����+���na��n����00(���6�;'ƾ+�@K[v�wS-�C����Y��q=���#Ǭ�Ğ����3�����OZ�R�gNΠp�_�&���P�P���o��`E�i�eBz�k:z�u�#Ԧ�����s�u긦#�3�em��`z��a1Z�G2�q6ȩp֦������r��0�<����Y��F�w�[���"0��X����,+i��{�F%�?��`[5�sr9;�����O��u�����5(��C��J�SkaAD�r~?�s<S��ټdY~'S�fS�
�tA#�M>��� ��	.Hb��p
]R�&A>k/�j2�F���dA��/�߾�k^��<N�\1c������B��L�M�*��u&��̭�2g�����>7�Q$��$y��lЪ˅�}F�����Ǽ�z��G�/�&X�Y�[��6x�1{s�����}ޮ�0	��>W��/rL��w ���|�c�5�I��w4ZBu���d+��3t��aQ���b�����*�z��Ԙ��[lU>&�I�(�8�{K�dٳ4��խG�� ����S��'V�x����%6�w{?��e��a8�%�<�Y/�<�%�Է��i]䲃��\��D�������z��mvƕ����g�+I��ں�ڧIS�U�(���������Vm����]G�)`O���OQvO뼍��-�TrA����� ����
iC����'bÉ����믨�vT�v�L<��7v���[jC,;���������g�l���ݢ���O��L���_4rL��B,��@PH�×�)0�}�b�p�;\F�7��w��m7qX�u������z<mGM�MND����+mM�`+H���d�3��<A|�y�g�,�g� ]�Χ	<�1)�I�c �h���|��擿��΅�.����s��B��O��~v3g:�˒�S�������-��-=�h�)lk����\T3h�m��i����_�7x��ks�\[�#����~�Q�=��4����Ruŵ��;���Ȋj� �rn�ŗP;�T*<O`�=a+�������r��ܼ ]c��{�f�\<��u�#��������ha�'.�*.i�)����gᅾ����N�4{ü��1��|�����<#bF��7��ѭX�l��:v�O�L�,���	j��n�J��Y�r���~��d�.@z�>���� �W2X�'T����� '�@���j�+���|12V��j���p����*�Ҫ�|�_+tx�\|Jw-�Nz��G�ހ��9��$4�N�LI���� ��hU���4N�I~�\��-j7�&�����~"����U��l�q�z"1)3�q���e	K���;��S��17S�#�I�$q:g���Υ�%�*�=�W��E@�-�F��z"?��x�;�G�"멹�/O�2���0�����Z7���������ۜ��d?y�O�x�X��c�`��=�W<k>��]N��|nbr�?��v	�^y8{.�ֲ3�/iaN?�.�s�Q(��4�5�6���>���d�KW�vW
�fi�9�/���D#�oʅ��M��	{�lؕpS?����6T���L3�	Y����w �#�I��H��;�D�Kv�_���Y�U���@� ��zE� !��NR�z�d���\:���=�Է4�<��������r��h� "\y~�
���Ť9�~��d�YPW�Vc�o�[�I��<5'��m�Uv��m���� \�7fA ���X;K��'���o�l)RO�d�N�Ws�S{��+�P����8[�� �$Z�����T[v}��mq�����t�ݸZ<M��YQU1���IG.�z*W�t�s���=���i!"���m0�X,,����a�,O�b9�z�a|�BV�%�������;*"���$򉈈"�f�d��ͧ��JH�����H��N�k'qRe�xN�a{� /�C�U�{�w���)R�PM�@H,�b�xpH�/��SZ^O��/Y��� ��yAD���e��&%�{��kBREw�vz�@p}@��k�J���`/��dH �&��\��)$�z�)>j�LG�' }�f�=�(U�`q���w�����6aN��XI�ٮb�J���[BM�;��b�$�Ts��,�Ͳ*�Y�VLa��URu�[�"x��KΥ;r��[+���N���A��}���&=C�AN���C�{I�G�^��˳��/��� ������i�..A��b��A��%- �/xƥ�������� �[��TZ-q�f#R�z�R;�_[��,z0���肺c=���!n8���߶l�R&��\kI�f��-u*�G�+�])��U��2�'�  �vRX^lt�����۸'��(�-�	憞�k��*םr��Z����=�*��ދ,�Ƭ@���M�����c��5�x�:���P�])��K��|
tʹu:���1�W�Q�A�ғY���jR��� �JPP���C�{g�[���K��=)��Um���g\���j���2
�	�8]������+,D֭�1T��ˈ���({�ǫ�hLFqr�f�e��%$�N �6�M7��1y837�z���+؟�&Sb� ��樫������f��!����C�'~W�_i�]O%�l�Ψ(�4��Qo�F ��P�s�|e*Nh:jų�@�u*6U�o���M�ZB�MG��vҗ��{����^��}F5��(�_j��n�`��Š�B���+��I�Y';��	 f��>rw��Ψsn��D�����7$�+�9�1�ҍ�1��z	RtEmV���jL����;ZΞi��W�A	,z]�U�l�苾n6Ou]�:[��6�9�@UX7'��ſD�Qh�� �&X�Vn;k�Y,�F>���H�������\�������W�4�7��5�c��@��U��G�`���t�Hx�"}"�$R.g�Ȓ�� ���_�5Ł������.-� !K��P	B��%f�h����J����5��%@xow���geemln� �<9����O����4l������X�6��(�����p�$�0��h��ǐa���\��3��a^� �}�_ȡY��}c�N�*qן��u2�7�?��g��(��x��*��&��V�M*�r4&",	]�և���[�%=���'�&��O�iV����Īyy5�
5UU��Up�79�ԮW���/�ԸNG���y@��ϟ<���Dq�Ν�cXqq��k5�:��x����`�?���e��H� ve�C���Ԥ'z��q7.�" �����+���2�����D-,|�0�B����-25�n�����͐�D�aXX��h"���<��!tr|�mؘ�j�
�B4�nn���|h�/uvv�Dt!�����;� �z�3y���4 �,��"j1S��|BB����r$��q?�=�y--"R�XX����#	����c����8�_(��P��g``��+q�G������6,�Ձ@��h�L_WR88������֟�M�ݤN ĸ����]gOG���GD �6�. 3���m����-T�-ֳ;��_AS�|`�Pae���;X*1��v�����X)�LP�5h��.�x�ID�I4�X}+¯ߑ�XbPXZ�f��F�|�M�n2jA���{��;vn_Y2�d��Wɰ D���]�ʎ�����6�����h��GAʛ�_f�C�	�^?d�z�������A�z�5U��'��E����}A�{�lY��(+�})��[�d$�^�j[X���8��h�g�$����e�.
0�O���S�M�A�����[��u(#�+�[a/2c/>�f��P/���2�
n��bt��B�-}�>�w��r��t����iY�k���F�M��?o�\BFZ�g�� �qhK}�rs0�<������T�(T�e�w��WW̊!+V�/Pd6I��o9$)2�N��!�^v��?���Wύ�}c`��$d�!H��	y8����M�9�;��j�${��,Z</6d��AW����I�#�1����eYe���ǭ1�k�C
���?J^t�z2$��}���V.�ug�=
���'�,?j4:ho�
2ē�ojEO��a��.���!B��c-�*���G��Ԯ�SX�Y���3�}(Ґ6�����U)�H?���;qCG��" ��<��3.7m�`'"^y�2 Su�	�Lf�=�8�i#�j#I3�D�/�wq��s��m�A��N�@bL�R��Ҿ�bP��>�\��|'�;*����lM�2`�m�P2�щ�<16�����l�0��jw5y�k�ĭK0�2�fN�s�m&���)���65?��-��!�/�1L������H�L�J�=��Ӵ9�4�E�W���}�zūM_B�
��.�"�Y�X?4�:qM7�<�9�Qp$=�mp�nn�����LҜp��s��>����b�2S�^$߰*Yt�4��ݰ*�R���
�� ���I��4�d'\����P^jhr��l����Gq!y`���|,m׀�xIb��
��ٶ[$�ym�X��^ۂn���ޭZ�A>U����Ȁ:�+0��1�����
���x�ה��:/���jav���V?�����=�SN&L-֥佩��Uz��u[�s�����3,1U�dEi,�����v�q����a�K����]LS2�N+��4s�A�������<G�����PgF-onyܩ���;XN}�җX*E�� "��B�A�#ے�a��s�AWS�	��&Ig����j;���]{>x6�'�r�^�qy&�;���B]�����UVs箓V�F����+����>B��K�����_9Y��8�gy�-D�W��g�ӱx0��o2 �גp ~7��h�qY_1�'�:��ܱj���Zo&�>�A1苈�"����.�i�f8���'���n@Mj:��OS2�����%��Ƨ�Ȭ����}����x��%[��Ƒ�PA�O ��$��x �W.чu�������|D/Sp��/���-���
儃�؅��K
F��3���[$J5�c�_���R����f}�H�u�;_�O�T鞴8����Z��;���Y5z�	+d�O�6 8�K�?F�_�e��r�ǾX�25TP��G�r�}�x�;( �>)�`/#D5D�o=;|��SH��H�x����贠�$�.��U�v�^?�x�1
����_�Ƹ/>@pa�d�|��v��I+�Tc�$���|x�cJ���e��V8�듗����n���Z�fE蛁p�iy{����9zLȞa1y����t��Z���Vm�K	�gPXk
��o�{�)z˧��$�j�š;2�R0�ʃT�R,N#�z���G���E�{[j�ՙLҼu�ϩW�V�h&[��� Wbb�zO��yy�|c3��CM����w���>�0���.�j^QqIO�U'@n/���f������x���wI��k0�8�x��^MZ��P8��$$?���_;ު�m�|���m	5�Z�M;Y2��&
�{+ϫg1�a/? Vb��l��)�K5����8�5w�@kc둈x�q��{�礼x}x��i��� aJ��n���v��������y�e6�1�;�u�Q^��̅$nt�|�s��E��������0B-'.$A�BEv�S80�GVE�؆�El�A�F%������r�r�*����m���� �ܢ���O��BV٦�F0V��<
���Ԫp<#�vI#�+��(�����הث�9���߱H`�cU0H j��a4f>�K9���5�oc�{����.n�Il.T�g̈ϔ�W�"�%2ֿ�U�����S���rY��GJ� ��I{�lq��o�#F���rô^���zxZ {�%u/V&v��Eb��*�	���U%Ģ~��j�v��~�J�{�G�I�\˦ڻ$L:=��δa��bW�D|ڷ��|�����sk�L��c(��=�TB_�/.����d���wλ�ᤧq�Їt�J#7��)��K�J�#�p49�2;��X.�x��:1���f̈́�*�q��	�wY���?�&$wqO���v��M}�	�ZiSmv���{�ބ�2?. R,��1��� ��,�yB�%W�x�7ܧ�������(s�7�B�F-�>�(�i&�Y�t� �I&F
@xJBx��wsq�~a�[�&���$�Q�}ɤ�(���oD�f������� Ā
|������k��>?i�	4ɾۙ�>*^[+\d���͜3��Ǫ�}W�j� ��ӭNI���@������F��H��8��$\3�z}h2��7�kf~�o�^>=��zs��+�F�gԻn/��Dc�_��kMԯ���}���s[C|1�[�T@:��
7���E~�ͯ�{E}��-^����Fm��ClQx�(���U�Xz��V�
��|�f�Vj�Oy<�����Qt��y�r�D/}j� w�!Q�Ldy?���7�:���d �RKp�mTr��e7�t�ov�|=BT�J��frN���-���
C��o�M���i;�J�C�ba��P���i���C��Ɗ}#�E�
�����d������[�%v��X	ٕ��|RX�8�E{�Nȸ��ӽp��#����a����8��+�\����k�\�I{Z�qc�C�i���>Μe�\+D+h>�|�Q����N��[E5�fa�����l�1�� H���h��%�U��U�y�hR���R�6r�I�J�6��Ƥ�
*N��ɲ�5j"�lArs�iـ�P���m)/��>7�nOq�,�m5Z1�oZ.�X����ͲkUYA�^���A�?�tX�x�����n�:z?O54!�aQ�P���k�Rgʫ�����c�rYV�U}$���e'O9'�x��g�>t`����MN�c�p�ca�{uL��z�z����2�%H�ǀ�v:)�a��,��(�l���`��l���xq��ag!#G�y���t.�ߝ�W1��}U�#����Q�I̋���C�.�Օ�;����E׽dX����H� �ܦ�T�3K�?ݲ�pm�1<��]y������ ��7��X��\�`�f�n
���t�k��^�o�%�<)���h�§G-�Mn 2�&����Tk�U&�A����mɥ-W]�����&��X�Ӊ�����=GU���o��ss}�e�� !)���|��wN�^�X��}CZ�O�eJ4�J��gs*���S3?��"�ƿ4]Zp�e�V��c�$���RB?������f��O.�yc�3�"\��?�?�.�a���ԋ	���7�qS:O�J�~DU�y�-;�i���ʓ��F�*��J���I�j�2�����QQX���rz!QC�F��ט��./�-<�.WP�Q^>�pN֗��?+�u6�|���e����΄��b�˥W�A�з����U��g�>q�^�`t޿�80�Y�0�Ƣ�6Ђ�c*�_Q���_Gd٧=�V�U��(7�u"���C5u���Vx��;@,Ǜ�@pa�M���p� ���J*4��'�r�7�3������>�x5λ�����Zޤv����ǿ��OJص�y
���ds�w'kn��Wj�^��I3*�%BL|ς�-��-S��/Js+cBP�z˓9��7��[=��+�s΍~����~��l}QM��>ӫ��>��'z}��w�H��
�/��W{f+����;"��&Q��~�L�I5���B��S��y��J�<[	��'�.eAUV;sՊ�&sF�\ZLqx!��|G�q
�����'޳�
��CW6�՟��  �x JE�<�>�z2:x�|ٱ�<%�gx5���g?�X#���&`A=�Q�Q��c��FJ�4:ڕogR�Hp���og�z/W����նÔ�V��:������ɗ-�\V�m֥<���Uo���[��(���6���7 w�EQ{��&L3F�ӴZ��+�@�Tw��h��x`�+��y�̚��o	�� z[�i�U�'��+�z��Hb���{�D��9.�֩:J��Fh�h�T�V�3Y7�	��m{��y��!���/��m�ǿ�:�T�ű(j��L�#� ����{��o]J�II�Q���{ɧ�^%��O�!YW8֟�y����L���8v|��!��.���lp�R��[Ɇ�����%�@�j���̓��ӸS��z
�^}��r���c�7�L@�����M8�l�)�s(�;!��QI�Ƴ0p�e�=��Uu 
��|�zjVx�/���"�������T U�,�N�umf�O9NC:VE?�T����0�.�`J�w4ZQ��3��j^P��k����ysl[�.,��S��R��J�60L2����70�Gsdt��<h��ҡe�m����$]΂4��y�ܿbUû�u��?w�!� ZDj���ۿL��qX8E����L��2>Jߤv]y�)��\_��� �����뮴s���ۓ_�&l��J���|&w��%�u^������'�^�Ԭ'GUN�h.V���l������������p�,�kJ����yi �W1�_"Y�a��RÞ[*z��R��b+��#@4��r��|���l �x�Rg����B?E<u�,&��Z�B��ە�ۛ.0�x�F����Lp!����KL����[b�<C�M3`���v'��Y{u n��vG���.�<���)R�_=NK�T�
v�XRx�]�r��p9���yz�H�2���~��R��k+䝂��Z�mb&��!>�A�����LѢ�����25饸�$�3��NVk�O��Lb�ЮΈ�k$��k�����$�ڞ�m���J�Eݣ�c��z9�<[;�Yd����
XS�/؅�d�S�:<n�_�����`�1րѰͣ�^Q�0�
�
��-�Ё̡��^�<8  �g�}tܧ�y.b�s���e�!��G�����6�͂��ں��pA��	����Os�P.���W�q,i�pY���W�`zE��^<�y/��d;��Q�R����@aɴ���I���x��B d��ϭC�ʌ�޹=iѳ��]�k�k�k�6�Y{��@Efj8�3�y�B��޲���ݶ�_��<$�L�wSm���X-����Y�d5�yƈ������ϣQ��ϴD�6�����4����G�JҖ�u�W�t�!����[\;�C�(��V�"ZS��*3e�����=�5��d��^�l\� i.�5wLY���wq�+o\!rg��k�I�R��;];�z�`p�eF�-JZM觬P����4�^/2�~03,�EӍ��lq�V=��7K���4�Z����b�X/�Z]|L��w��r�G�Wc�@�����A�H�;�?��>��O>/�/v8���R&��B Jt�~zQ�7�f����*	��r��I:=��S�s1<2�c��%�'CTe���&KMkq�ᡦcd����Y�/ٱ/�v��N PN���HD�)���Q�*a��������H�粱gP�Ԍ�⾈GN�Jb��ij���"i�9�z�eX�h�2^%L�1��Ez���N�=j�P�ɘC�P�J$y�� �u��n~Am�����ٍ er���0�:K���h�8��9 �,T�ֱ��5�P:��or�}}%)��z
 ��:��<�W�hc�,�;,���a�Y|�n��:^ǯ���O29'�ܽQ�����+�U�,T�29�j��&��u��_z��q�7�W���������]Em�R��	�p��Y?&��wP���ʩ�U��� ������vm��V�U��)�l�/�� )/Gk��k�;����;���wg�5AA
�]EFf�ˏ�T�n�`�B�q�G�G�F%Cy��RDj���~�b��ID�"�v��6$�U��X��wD����2��<�� �x��P�].�
;�Q�Hg�����w�gy��p�ӭ�e�h9��2��wY�o	{B����� ��.� �Г�ԛ�V��� *ռ}A��L���QmX�d���n�WI�[K�*y��b�Q����/�B���Z�Km~�ف�_h��R	��c+���+²��V��)���9{�������X�=F���@�p�r�[��
����Aj�W^X�C���A�-��a�M�\u�ZrJr{���������Zz]����u��\b�v��X�Y�o��V��ݛXDN���&��y�֟Ќ]=e�)���p�f��8	��Ŀ�:�;�9���&��Y�7Q��ܥWϥ#y<^Sg�/�'��D&��vUs�*������Z�<4kn�Dկ�5\p軸Rѻ??D�hI�G1���mD��:5[@c�Xo�d}��s�$�k=!8�Հ���-M}�a,�nu�>C(J'��Riu��L]���;+vazkd�	Y�P�,E �fҦ�nbR����AU���#�����5��:Z�џ��ށ����v.>�tP�oF�N}��7oi}��+aiJ滔��?�o�Znމ-2N�B�D�@�� ����!T�G�E�f`�l�r
3~G�,��zߡ�Ie�
9$���c*k����Q�No�,�*CGhW���͵q�7TQƷu��IrΣ�vUQ���G�In:���)\������-�xD�Q���d%+8K�P��b�J #й�%�w8�6���˽.���җ�Y��j�)K 2qVm�>��E�YF��u[��)^ܝ�P�	R��{��R�����ݡh�C)P�]��[������A�Y{�9���&���d;�E�vZO�2�nGE��������D�:f�!���b��Nt����M�d1�^�,��G�X�5�3��~ٜ>Qq%���e����Ѹv�?E!kIM��Ii�Ԙ��D��n����n[��V�j����u���r��~絓?2rbs����_�Km�Z�^���"�dS�s	��D�_��#�6>��y7���=LG*n���4Ii�8��N\
���������p�@�-���,��[ �O����	c��Ij-�FMZ
�`Z��m��b��Y/P�d����gǻr�I���G��z���b�ߙ`}�����;+�?�`�F���Fk�Ew���P�U~��m֬�@UU�����GA�)m%�D�-��\���W7X�{\0�m�2�(3Dd^�����(V�M�#�����@�#�=[]��'��#N�;���K�>!;��3:����;��xx�LL��	�#$�|�L`��mQ�F�d�M$�%�Zih.6Z����MF���	���?:���D�]Č�)i�B��4���T�d(���qb*Ktt��p}��}
[<�7�N����_-��d)S���{��������f^�\o��&����v!C�F_�#p�@
�1�s@�xFL©p�)5�����v�";��(���z�&ϙr���j'P�^�>��1��'�ϳ��{1ԯ� ւ#QO{(���}B�~>ߜr�'����r���^(���W*�p,)����	bGH�U���c0���;d�l��<qּ�u��/�d?�r��7�˩���h�u6���I��v��aWEBBN�YD���q��8�Ua�R4_�Pd�1��4�^~iQ:�в��]F��S��Ͼ���\
�{s����UT��?0ܧ�&���3�d\m�+be.�[;��W��/I��@�eȓ��r����:ē�F ����Ԯ�m.����6��3����~���ۘZ+��=�Q́_�^.��He�i0����z�/X����?"�>�Q�U'd�0���f����ٲU_���ÍLq�v��w�|Jq����3��8���! 4�y]*�'��b	Vzn��=�qN�j26>m/�x$ Ňq���UWv
2��<�i��9PYu��0��w��W���U�"%�l�i�"W�i<���q�Ԁ,
�E�yVM���C�������k`?��oj���n7s</~�&i�Y�0z��^���#=x9��m7628_d��*�J��V�Zu�ҏT!��X���,K��d�LW�S��[���lً�4)�-k��WANt��%�3<�힎��s(��O<dZ�w�GG�{6�]({}� ���O#L���$�}���p�Z�\]�e���"	�!n���T����G���@F�\L�Ҋ2���msA�N]�#����&�I�C�"�Dq�?����7K���gA8��{=�b��C����Y!�?H�7>>Mb�@����kq�f��k�%<O�v��{��|�?_��h�͛�=/[��n�F��`+��;7�:�h��Gtl'l�n�3c�~�b�\aG?ݡ�����s��:�ԧ�5D���F�\�G5^�Ӡ�.ӧ���.���C� ��	v�	�(�:k��nT\���D&zX_�{*l}���Ȃ�&����8��S�ߏ	r�r�e��%+���@��w�
b�Q!���g���r�������}B|�Q����L�}J����/��J�ec�>2�rS�3:�gޯ��|��B���)��8ݕ���h��e���_6�
��2�w�\ t�����z�	�.�-3�F�(h��b���q�p��t�s�>�خc�oF�!�����j��j>��R���ҟ�6�k�b��v㬖>����Ӄr�_*/�}��f^v��M9��7�@(</6��]��6�����0=�~��o��WT*�~�|�3:_�z�)���c'��Em}�@�sd��e3:��q���2W��A)��aB6O��Q�J�����C�O;��{��L�:r��ڽy��l&E�����#���IaA5<@]��kn~��:�b����}�Q�H���ʊ�p��I4.� �c�7��
���@�r�7�r�d���<?�ߧ��?������|���E�Sxv;�]�AR�}Gf<i&P��c:P���j<�V�	v���#�-�� <�� 1J�[��;�����4�A!bj����4�ũ	�̘KN-ʼy6�[���ٓ>\�r��aqѓ�b���a�'��5�񥋚�z�)\��/�؋���	�zC��>�|�������E��E�٨��s�|I#\�V�Uf�e�^.,��f0����ׅ��q9�}� h�2�uJ����=�*(�z���\��X��K�5˙Q��*�߆B�����jǣ����2CDPv����<������b������7���T�ҹO;�j��eSl��QE�"�R�*fKz^������� wj���}q\�l��R��{ӑ�n/���U��#��,l
����I�M�Q��8�9���H�ͣl�~h`{�S�>��X�V���85��^f��M\)1](��^gF���:3Y)�@�(#�����z������cy/T����k~$ |�wnx R\�P���i��%����	���SA�GR)ȕ����P�u�����F}	����x��gsT�s�%t�CH:Dp����.��(�uϮ������p8F(��~s�9�A�@�R�PRv�y�9ހ ;�K�)g����3���NA���5 6���~bߤu0��L���1�"�?����ُ��C�洼�"�1���PX�x����t�3��1��挣�Ͷ~�g<�b�8���rvȗ�S����2���Fmy�S��%Ty��P�z�r����r���z�����e�Ue�Q���� U-#����e-K������m�(�X��}�Q������\M ��:"!��*�j&0��.
e�FDҾ��٧����aB�pq��vo�
�O-����le=�&l���e�IU���kia^Y`��T1dj�|[�70��L�25Im1�p���ecەЗ+�~�;�A���5Vx*���œ�V�cZa\����䧈����\L�ԝSv��o��W��9{j騝�Ͱ[������"ɹb�=�
���z�IS�$fX�b2�@U^vi�Gvw2h�]�4GA�oڜ��ߦ����,�4���xk�%�@+���uC`sb����RB�r��pr}E�sZ����n&��z�ܓἦ&J�Y�������ᝲ��rM�;zZ�@�%y͵{��ȸ�C]��ݱ���������Lw�$�'�d��혂?�0�u�� ߉cI�]���N�3�ZGv��5a�"��F���[�<��}��A�m����z�_9"$�J�~(�d���s2v�Ȑ��d�PQ�	\�dH�:u��^�\�kjTTk n=�`y����9}�����#�|��}(U_���!���l���cb��Y/�(o� ��V�4�"*���V�?݋X��p�?� CU1�}dͰ7чd5V4��Z���#Zp�P��O�*��ޔ�_P���X�1v&��� ⶖ����d
�;{�{C[����Q�SA����J<�a���J�K���mţ"���0���Tp���+7SI���|��tb|Q�g,0z,�V�k����`���< w%>贴h���W��;R��K�ז���O��C���	���=���a�x~�L��뀮��m����r�+��F'�U�oE���61EψJ�=̀Xex�0��պ�a���̙O�)��ښ�1^�E�M(]�E�_^0�o�8~�B>���@���pp;��e	����s$r �x�x�q�%F�zh����?c7�|婉��~~fB��dP���I[�.n��U�|�<u��p{��8�SӇ�/���Z��j�O�J��5��F�u���}����!DK��O��>4�/�yK�P�	�b</=}qH6[�Y�h����ͭfa �a\��8�a��gO7f��?N��þ8k��$�o��?�B���_��8ۻ~��S\t++�J�g*u�吳��P����z�$ %��%�'U��/�]ի-�E9�k�u�՞�3���iM��~�p�K�`%35���F]�S��ow��	<�ԑ"���I;���M��v�o5�v��U�	���S�܋�A��mp���F[��fx֭�@���' O��F�K�.������,)rm�nx�Ϙ|�;x�����|���+����z������x����Oh���ʩ"�0��_nDIѽ�"@{>�ǰ��é=���2���PƢ1���+wƄ2@���5�#�+H�Y���|�g���0ѡ��٪3� �Z��u��?2[2NP�d��D�^����L�_�y�zT��Oŉ%p��~@��w�޾�I��3Uh�4��I�nS J��� ha<���t�|rr��#��u�2�kHli��O�Ʒ�%����j4�Y)������S��35K�ż��pȋ��u��}aۻ���<a�7��ţ�/�׹k�x��v�˲ {{�g����:l<�l$vm�X�j�U�M��8DR�j��yє�(C3�#ٲ�fR�m�aR��/q �7$�܀6x\�J�̘�A�|��hHC�/Ԉl�bO�o�Y�v���ƝM�J��{�b�)������l�+��]Բ*�~R3y����������ٯ�rj%�L:�(�},��C�lo!��Z�i��2�9Ny2;��ו	0}����/W݉FU\'�	��j �>�_r]��������OJ�6�Lx���PV�JEo�����Y��%��[9��
�@����r�
���&h���O�J�a���+H�գ�2�-*+�kk��0c�4��E諮ث�~K�0ݔW��G��D�L�Ɗ*��n
��F�:�v����^
?��x�q�)pB�N�<��CxU�a ��ME]
&���@�EX�Y�����7�+���?g	�@كt��ˇ�(�^��*�>v�a��^+xD�����hdߧw�<�N�np��J�#��{��J�5އ3�/>_�&Z{��a��m��-8��U��F���i�P�%�.agK'X�������FƬZ!&���_�4߹L���s��JPˢ��'�2.E����fA<��$p��ȉ�_ɐ��R��^Ԍ��4@;�6T�~@a(99á�˛
��χ*Gf,�c�!��ȭDy��^(�~q��f�A��2�yG�[��#
�k�}�T�y�whV�����`�߹!;4������e�*�na�<6w,ױÚ�2�˃�!]�!�ƛ�������F]ƺ��� (�_(E����#���ZA&�u�Je���`OHLf*��.X�'ad|������=�� ӂ��3JH>{e�ek���̖��:�Lz�4�qv$9o��tggg�_����b	�E�"$Ӳ�w0s�El�7����i1��<���G̯��1�ڜx���"�L��s���)�m~e��=�ʒ��uN����+���Q;n����#a%��ѐ��Sɗ����g#��J��"���9���T�Qɲ
��E����H�Է�꼘�$�?~�t"���������c�d�~ö��|`"�.w�V2�k^�>�����O��ԟE�Q"H8�2p��\	��M��3�a�Q~F�`ΰ�
A9	�(G�Y;i�L�h�R��?�df�|�֟��@U�k�4�ȘuO�s��j-������ ���C�����,���y
���fQf��M��D�nUm�w���n�Wx1�Um���ӝ]x���m�G3��5
߯��
#��j��,��+��*}�Ѓs}��ZH�����5��3�+��w���r���ƺ�]�-n��;YY���Q0�5�@������"�/S�G��
�݀J?t*f����=�Y����~Ѹ�G�ї�㆛]��1�v�W|]�����[�����Bw\���H_#�ƭ��K�}�˖�%ʖhP��0�y[��۶=�#M@a��t���M������R�Λ�!���&PӚ�l�M���tUp(��N4y���[c�J}O�dk\�x$�>�LGq�8�5����D����Q�o��6Z�xL�:��Ȅ
�l�,���:rB���='$]�E��n�W���8�$/�q��.;��?;������W/��j�q��!����󺭰,����LP�W��5����6*�IH��4�I��&h�M}x@K�@Zl�/�lu��Qi���е����tΣ��c�*��@����DI����zG�7�GU>:����Tu�Ͳ�m]F�������6>į�����xF2�ܓt�7��-)��=(Z)k�H
��*�W�,1s��>I����7x�6G�ME�b8�Yt�t��8��2��@����Y�_'`>�JG7�k��se�����ǃ�i����ϝK�D4�#b����t�����z�|W�X:�Q]�!VO&�n����V��%��~���3��z;sA��
�4�?�tmWRDEc�ؼ���49J�@��G���l�m��x2g�a�k�[ͫ�����G�h?��=ׯxO=��c��5�y;�h��,�N�����rAS{_��2I�3�v�6[٘;�Kd�ۣ��լ���6²Z֤�e�WGG2�G�ɺ��<S;~R~|-�����z�+��ٔo��Dol3G�f��C��N2��v�m�G,n~o�K��!MM_�2��O���7EkTO_�[� �����M�SdE�8BSit����Pkɹ���9�"��o��L���C�u+tG�xB�^�!�0h�q�B�0%}4K���<��bG����2��M,������t(̛�.����Hj	1r;P&ɖ�9}��WcG$`w�z��W��l?����*�_�ċ)��U���H��(3?%�2vLy��wt��$M�fd������d��܃Z\��h����IĘ3TjHʄ���H1,�(aMڪ���V���Q������+�G�j��5(q�7�v�j���"�@�P�D����BP�����X��Q�'GG��4e g��o�w�э���{yB��� ��X*���P庩�r��甑�;$�^��?;kڷk�2�]�~sh�e����L����R��1�DFއ�ۿ��Q�� 
�Q���t�A�7ub��SIDr����턪�S"U	���8�-+��k�V�o��b}���?DJ��n�L���KC'���#; �H*�2�L�oq'�I�]�ƺ���c��֨��J&P�<Ro��\bp���&��簿�6P-wD{������S��wXo���gh!2����D8�Z�P��թ�~����O�p:��Ω�iB�+���_%��<[�A�����w�����?R�K�l��8CN�����}\�ed�A�z{�| B~~S�B�����Х��R�k^����սt�����1���a!�|H�_�KԀKTb̯W��##����x*����x7]�,I�<9�nF���D�4����2�t��r�2�o��fK7�4���z6?�s���FC̝E!��U��]�M�-)|}���E��ɘ�`�'��b��g��>6���#�w-��S��r}%�落���<Z���߲}z+�9�5�p�>ʒ�#�p�kk4m�e��*������X;e�#d՛ ޮK������xt�v�����SW.tG����B��m���~\f���PEŊ���x`܋\fř>�|D�u��������|$���~�a�Rf�nQ��Z�h��Ǥ�p<��˺�+����ѹ��G)��n.:�h��,�&�d�3��ƚ�7H]���RJ����F��j̒v��M��B㽤r��';Q�H�>;)ސ�pCEpE�� 78���-�Ы��U����g�|	���8G��03��'��v���/�1/�̗�ٕ���-�3��L�B�Es�2�O���t3ｽ��I�c�Mգ?q�˴�/4h_��Y�)�U��Z��(z�s$e��w]�p�)�V��L��Wo�ɦ-q��T>n)#]�L����|>�h5�dT��L�z����� �AV���;;X��Vn�/����]PPj��
}��)���iF��l�(HQ�VkNJu��L������5$���� -�}\ium'c�q�D_���z��LL�r�R�e��@�(T�,��V#��c�k��0�5�2�v�d/�1㝈y�y��l���\.�Ks����ծmm�-R�<��$5�)�����"8�/�r�kM'b���JWyBG�h�0��s�P0��HMZ��l!��Ѱ�^��oe�� �0:��^���%�V�6���4a�|LП��J���9��u2�b~w�(�l�]�5r�%��A���ô���,�@GY$�Q��zlqM��(�:51m�$Nl�lf~��@oRƅ��IU�F9��wa�F�k�x�8��A�y�ݵ�c����G���Ҟ>R��z(�e�6U)�	o�玒F��$�Qf��V^0�+N��ǓGq�Պ񆱎��2ƥٳ'>0�^{Pa�_��31C�>��_ [�W0�\����oD��{�����9�?Ľ��WR՟|��U�����(K�����'W�}y���dz����)�{m�����;�trn��t\�����Y�Z�V�ҕ%���B.cAO����Y��}d�&�c���aP�g��x�>��_g5pR$ޟRa_�Qh�J��NG�Wܟ�ϮZW>���6�T��N	L�0ɉ4���sf�[j:��͘RT4�O��&�P>g�i&C�\�[`;5��$�s�'r�����&L�ْ���4�Ⴗ������ƼNB�x����+z����V���$B����C���eіu{��߻�䅭,��;�ВY}/3Ys�]Tf+#�� C �y)a\�(� ���T+�
Iϑ�T;6�L���$�}D������<"|�NbG�-�H���dTxj2��K��т:W� ��
2 m���xx�K�h�͹X$c����m(��K�h.*��F�fu�������5�x5�R%5�DD{	(C�#˲k`e�Hޫ�F+��!�\��\!���
?�L��)l��x���_d�>��<����{��,��&Zc�<���m��I�w|��k	O����!�Bx`]�O��-P�'�sSP/�:�4�!�wA�Z��)C�����;��Vu7	Ώp��@j��ҷ�:�9\#�Wi�8%\���=���0.B��"��:�D��A�8Ԓ.�	r\���/��I~�2ᤸ�MG"�|�@CHʼ�dӶ���Q>�߮*[�U�Lź��\v&�wsL�z��U����5�|b��eL�[��;x~Y9FC�	أ�V��A�̍?�l�����I�Δ�4tC��$ʪC�.�>��H�f;�P�aM�nK9oz�$[)�X�e�ˠ	Ee����{�|�]'��LAc��-�Ӿ��By��=�z��9w8RyГnO{-Ą*��b�,�N�o�Pw~��m�F����|�y��Z*In���YR�n?���{����x����BL�hn���U,�ʘb;���Az#��t�9����XY��&����?�t����F�d�&@[Y���^�NC8�w�Y쩭�Wʼ)_#��S�Y��V~'7���p���8��|R�>�����!�]�i\�G��3���(�7�����9���|��&F�jve���O�43��0���hu�Xqc3�����f�u��w,Uu�b�1l{7q�%�v����i'�hd��=Q4t�Ü[ݒE�Kz��0���az�yU.���wc�?���aJ��ef'k��l��"OT�	����D]�GKk�D:�į�_S�J&Z���:C'�L������|���#�
*������X�)SsC�F!ʖ6�� x��-�h������L�j�H黨q���h��-�+��sW�ڭ��{
*��c1����%r��9�ax�!َ��M�֛q,�+�1��7�==��^Lqˢ^F�P�/^}X@�n
=)���c��؉MhQ�|�%m6�C~� sx٬��}*���S��I��P�y�����u`_�^mZ��,ԔV �ʌ��E�>���k�3z>����$�y,kk[��ʏ�)�B�u�A�U���T2�e�2S<����Ԡ���fx�Uqet:Yd�cg�hc"Q�����t�/�ma"���.�<0�M7D��:RAO��@f�w£w���ª2�3ڻ0Iۂ	r��`"~=ʢ��R�,�d�;,��쭄�����Q>�􄶵�wUz\]�8pH����}�A�W;P�UԻ���w%Q"�����P(=d���������y����1�[����y���d�V�������D�>����^�}P�t���Jm�n
0V��|�]�;�F��I��K+�ºFF���<�Lz���7@�O}�^:v	3h/^�;H�K��`�5�2 �������t�>�C}~K-��!�A=�?�z������h��AR��V}�N����ל߮���x�|����0�� �Aw��j2��C��nuߞ��}��Kz�A1kGK����JiU����w������]�twӷ�(�~�����0�����k������Q ��$G�:U�0S��������w��}����~���ѿ�(��YEk�qIѡ�!��49#W]�<r��:3��'�����z�g?���[�/}�Q�ؠ���d#����P�#�`�ErD`���}�*�K�GN�
/�J��P�6_�u�ld���Ԉ�mA��M��SQ�}~t�][�h�a��F��y,�	��P:�0*��E5�8��䔨�����t��^�I�_��k�G
Nh�뉀B�{WPG�"�i@�,��ٍB�-砦6u��7��|�T��a�����N\�ø�*h�l��7>'A�i<��u�-~6�B��Q('��w����O�r�����qI��X-��U�3�.�������%�n�a�1�1� *a0��K���va>�����ɱ%;ɫǝ�f;��kZ�����BA/�/9���J����i��O7 �B����BS[���w�V�v�b�?dJ��YV����`>��c\������h��z"�
���%���a�c����4�d5T�o�g�{���|���t�;���@�k���жA� ҍ���ݟx�HW�8�F��"GD�B���h]f\S���3���
��(��5P �O09J����	ݣ��(��z�&�T7wϲn����$���N(���~ ����~&��OX�#�4m�t�$��]f���.g�e2�m�����:$7>l��Z���1���#F�M�#���ɝ��Xa>?5aw��5�/��Dy�躙�ߣ���l[懙��o��j��|f��{퍼�m� ���<q^~<�](�R>�2>b"؝�O$\��q��U����bد���J֡p���g�=�zG�^��/����Mu�e��B�`��h3�[�ְW�#��N3�Ω�9�rֽװ�� >].Zz�����O�0�۝��:!聀u¡ר����A�X�3l���3���_݆��7�d#�D�_�*�6�>�)d'��(�k0D�qǚ6(;�(��\\ֳ�Τ��"��Ѭ�h)�i ]��� ?Goq�����l�A@o���|�!7Y��bm�7=��NP��Y0B�5�p12�Օ��:oq�R
�,xi�z�����Q��4�����ޑE�W�mX�v� ��tKA�����N�Hp*�$a9�j�}uf
2m2dv͛�,�"��H���4���o~�T�싶B~�!��>�{�^��u�',�Ď�΢6qd���M�1��5#�������l�ѣ[���%��񄰀��t5��o�{}��|,�J!�=�_�bE�#NR?���D�y��{g1哭��-
�څ��*�6V�73�m!��du�;oz���W2����j�/'�r6,o�8:� KP8�o-���t��P/b=�k^��iQo�g$Wsڸ�=�z���=��� V��X�R۪�(|����Û��bo@�5K�s$�P��:��q�����Y55 >w-a��.Ub�0���\F+���Sد��� ^B~�lպǺ诓Vԉ����(�ff��uh�R�@v�34b0�!�%���)="xpF��b��B�7�POcg
 @�lՉB�Ɏаx��y�Oу｜����-O�4{�}JeXH����naK,�� ���\���T1���j�)����L���r�m	� �@Vo�i������ע�ۓp9�j�Y�<�du#g,��A�2y>��ԁw����L���ie�k�&����P�����@�-J)4�r�������@2�_%�5�����Z��8HK;$�T��3�M�����Ą��O�"������r&W��s���c�?  ��!���R���9 =�%'3�֤���o��v�F?� �zx�-m��u��p��s�(�8�X��4���xd˹��D[]�b�#TC�ǨjSAǄ�\�Q����g�>�gĻ�9���o>�^��E�E�E��g���z�3�_l�b��
��%�Fw����C�n-�1E�`�%������j@��6�D���F7)[m��)�}J?
FW���%ܢC d\�"H����@a&I�&s�2у�N~nw%ʖ�r\X%��v<������q�(�c�����e�`m���f���0O�n"����Vhu�^c�=��j�w����Uxr���_�D�f	��V�I��w����V%F8���]��1����?�s+^Qo�������/+:'z�辴 �KޟyLu�.A�2�|GR��������j%U��V���DlG�㑛X����Z��ۏ.��M}'�_�$و��YS������;%��?�q��!	����U���'���������3Ͼ���U�bLN-�q�W�6Ayq�r�ŘҠ�r�T��=�p<�c�{�۵�6򅇩7f� |P���n�Tf`#k9�R���3|�Ϊ�lu��Aa���$<���fE�Q�(�C�"ODv^�"��cH1��r�fl/
y���1��Q�Ҟ�g��� P��\�t�!:(1ڍ�&���T��3�M�<���~^|n`� ��n(��%�`��5���<?�궜��</��D<{�J�+�sa�L�{��g������% =�<�n���LװU������)ݹ����-bE������������Ǧ���+6J�[Ȏ�)��ȕ�z�M��h��4�jwv�'� q�ԟWwlw�6S@	��#DG��u}�L���0�:TDh�Y@�����lS4��CT���u� ��(�u�tR�\U(��^�+8����t��4�R�Q�!��J��.n-$�]�_Ʌ	g7z)m3�]�0�������l�n����u!Qd����}�������|������]��q`[v�Ԇ�P�{�V��Uo>B(J���˦��#�/]���M"��ѐ����ikj�Y\�N=^	O�^S���y��VOa���؈��`O�Q���i����E:+����������}���V�b�H�O$��������,�[�yR����{���7�p�W>9}�\��S"��J�	�W�:ݢ�d ˨E4�s{�q�$F����D�n�K������/��_������<��у���+w�޷�J�|>ZĻ粠��n�A�����@�ѝ��±X'���ՙ����)�����.cAqGS.��h�8}i�J�8"�P��[Yd쉢�-}�y簙�ĝ�-/�(��0��=[��&:LZ�Ǽ�yH^ZW|n�AV	�����	+,�2&cP��qiņ�ӻ�S���É����}��yXU[�]׮Ʒv���N?���b�E�o�{�ctp����|g�ͽ9Hي���}3'�E .����b��lٛ���F�Xo$
�4�q�g��#&��r�������TyX�<�Q(`�Qn��&�Y}��'�$H3ĥd˃w�+ɁvoL�Q���0�pKoe��g�F�[̿j�]ʶ�D�-�K�[��c�K{,�?�h�>!�d�0?Yau=B,�����/��<����/���Vle�_fG�7%j�:��ST�8A'����/]�uYeN
�;Z@'ⱻa��Y��ص��������3M��nwsM�Lؑ�$����v�g�f�ϟQC�q
�g2����̞�����&��?�p̓�dŢm"��烫)߫�a��}�uu�r,]���ZŊ�m�kmz��~����m��'�����y� n�:
߀����̳���^�G��8[Wr���'�D.w4����K	�/{��/�cl�g����9���a!�����ͱ�P)Ѧ�/�_7#ؖ�E��
9�m�G"	��͘*{Cŏ5��,�0^��`\��T����o���a��Xk��kAp���S���xIX�볝�iU;
����+�+XMtnqq,���/��=��$�r�R`�����X�@�U'jX5���2�5'����+2'���|R��}W�=$����gF�2m�>>;^ 먨/	(�6d�t�����=�����#�2�J��4����d�x�?�@h4�}�o�y�M�����H��q��;��}��KX�N�<{�����܃T�adka�5 /�,��>;,����͍�?���[ɗ������eɨ���b�5����y����/����'#����з�����N<�:�J�̶�%I>giV3�O���Y Qt�J�؊��Io3�ُ�Ԍ�OH<�0�J6P�&|{�m�B�W!*S�G��G&��o��)�ZA���T]>d��G�Gm�Q<஥�l;j�m�3��w5�҆�_l����aj��,�ؓ��Y��)j��NM�Z�oɷ��H{YhT�������Ǆ3���A?�����3͌8�C�E��&�-�4��i[du�=,:��&ú���#��6&���d<�j;q�&F+���J��7x�����i̃�J"�j3����j�z��S5��j&X���Q��sS�JtW�)]�{����&�ۼZc��p�-�]J3n��w���p6�G�!�*�UQ��,s	zE��w�οQ��M�?ں
}�BK�F��#`�e���9����q6���"%V~��k6'��:��k֘�#r�,g�
Pk|ĉ��1J�"�ĔD��	�zߨߞ(�]��+8�7���O��p^)���*j*���2E����Z�)�Ϗ	��O"��<��jO�d�v^���|���J(�e�$��9�@��@Eod��(.}�R�/�wd+=7)��ǏO�O�{��G��&�=W�u�_y�l��J��O��p'L�����3=4����RF^}2�O���k�\��O�U�� �:��n"y���h��/12���|���O���}�Ůl�!c&������	Y�����⁥fo�᭜��uвt=-S�P����P�{�[�*����Խ�o�&�k��"^J,��ך�"���/�`�������֦Q�l�?�o�
6a�|F�]
+��'�X�i�]�m�k6�w<���g�+��:�o����!w�ĉ���L��������&��3֟�9d6�j[���n'���WL/�\'|���|��z|㽐������-K#��L�o1�1�P'��'ni� ��7�,���iy[qͶ2G���p�y��F11?�r�s}�%�|4��7ӯD��	��V��7��zl�V�'�ޝ�g��XZAm=ط��L�8C(̄\YV�;b#EBJ>N^��5��H��zA���V4<���Š��k�y�U���~���
FQ
�ù�eļ��l]�3ve7�Gͼ�ɍ�v���u:�&υ��#/��<�?kX��]��!����"2�(y~�	����.~j��3W�o-9��M����
2{Q��͏	�|���l�U���q�M#m�PԆ�?gdwWlbC	����7����%�?��: m�����)�O��4�F��ù���~o����A=ɚY�����"%v�d�g�.}¥��h�΀���4���AJh�v#]�!��;]!��&������.X��.޲�H[�2̲o���Ci��-O�D�3ō�M���M\��ML�Ɔ^p�h����YМ_��n��8���e�)Lw����~��$��9�B��Qt�z�?�E��XR��؁'�7��I[�~���ª%�4N��`T�f�0T]'��:j�ň9�v�ܞ��șB�����;�\��=��n�&�]p��[y��~�0s�_�-������Q�Q/�5JZZ��d_�^�+�����u��J�m�^�G��Z��W��:�g��D�ek��nOdF��Ւ��穹`�	�
��NuqZ�R��?�0�U_�g��n�~��	$������~���'�jՋ�,5b�L*S��������zc�a�ٚ�%95#y���vJ�J�Ď��:�s�;KZ�gb�yf�yo�A�|�v��72L��Dڪ��Ds�3���h�5��k���m�Ջx����IWe��_����6�Ek�<�K�z���zB��_Q3/��YS�OÉ�{\��<�G�W�ձ,]t��.!��Ɲ��	��A���nA�݂��o89������f�{���V�ջ4��O4�����m��I���9ZS��k0/�
 �y�C%��zj��%�>�Z�|��R��Q�	�в�ϟ���n#�kW��ܿqid�7�B'v��4�9�ENP���̓MS�'�x��Oh-��J1�h`���DJG�g�=�I���Ȅ��s]:��?Q~E�eR���Nt��)�n|vd|�{gd�Z�^����%��ݙ���50�D��a�i���ɲB翱�N�b_���gU�PU#��5�oJoq�4CW8�u��7���mK���u]&�h�*g��&&�-{���ùdl�4�g�pu��,_RI�OCea\�(tP��Z�+?<"��A驍[�2jW�z�J���0"�L��%!O�PZ[8�܅��۵�X���?5�r�hK����n��K�Px��3ǎ�1e�~0�s޷���م����[=��l S4�]��"�E٣�L�:,�E����:�/�:�0�+7zZi���nO>�H~��daH���/.繷����J�1,s6�rWǗ��@*��
]ٛ��R2R~Pn_�V
��ٱk�I*�QQ̺�#�)ClHY8���o�g�2�Ȇ_��˛ �q�;�� �	'�^��Q'�� ���t[,�����4���]m�(�~�ty��ވ�Ju��z���`�H���#��O���1�ұ61t�X2�E��6*.z���$an���U�T�b՟:����?�Z���� ����0m	���X��=��U��_�m�g~(to��d('\5Ta� ��	#N������U�j �������%
-��$���ƺ����y�����P�(#�(�mUt��<U����P����p��O<Q�+���P�V�?O���rɝ߀C<��5��'+��b�M���$��� �<c��c�a)v~E�ō�0��؛�AA�q0��g�����10S�a(Cz��C;��`;�4ý<�-��㎽9b���Y��W��>��*:X�yW~5\��%6h*F3;��͚���4T,��Q���(ƶx�L�M1�Mkr�tu�2aņ�Ucڈm}:C��0V|"P<�2��J /F('^���b~5EL^��v,u ��R��o��Dx:�`��0[xX:L�[P
�R<y?v��1�-�s��]>�}-�z��0c��&��O�q����`#0@^��7Oe�8�v�1[\��1 Ys��I~��<�N�i x�1R�w���Ucn֝Y�` p��y˖�ɝd�1�r�xP"TD#v�����~89H�	�Cj *"O_�`�U�,D��2�t��Ht�Lr擻����u�#XU�p��G��R�������ݽ&��<5H��W'8�^V6 /�����)-�CkG��
�0ɚ6�9j9�K�#N[�H��d�K<�?��BE��ĥk ���~xG����<H�eH^?OA�"����]8?_:�h\tB�ۦ�5�<{:Y��y~J�O�Jf���ƦOqa]bz��7���|�2�48�C��q�Ɍ�{Q�(i'a����ՙT���%��0�DHk���h���xu���O��!�vN6/W$��A2oX��	�z����9F/�5;ݻ�ڋ�T����)6�F�<��8��0�9|pN����͍,��3f�i!j�`���o�:����{�X�Ӊ�Z]�[�c�͟5��
#����JK�I��^X�}��Z|�`*��o��j�����Fyi/���y���rj���� M�#�Y�ӏ�_Q�U�;@[鶩�#��۾��|N�t�I	
�֒E" � �� 0yް�wU^�!A\e����O�|%��	K,A��=���#\]�aIK_���o�-ED�8�E�9/�������)T���(ı�:%p��i�V��.D�Z
��V9y�=e���P>���%��
�(H֛��Ya��~���u\*����=>	�c��"Vg�~��9.@`z�.|�Zu$�����A��ગK���p[��h���V� �����쇖E�W���q̻"���jn�E��jD/mH�ƴ�&H�~S!5`�+��{SO�F��kS����(��}��Du+d^c8}�b|\/�$^�PAd�,0�����t��1���=�%e��˷A��@C�1���[MF�u�tü�m �Y|�$
"�J,^��â�m��f�#� R��b�;�DQhT�7� ��h<���@��J�'�{�K2��>�F|��h�7ˎ��[��p�힖�8�2Vn�X�<���K��D1W_ѫ�=��2>�Fӈ!f�{�T=s�SWg_|3�V�WSbn͎�<$Ù4 x�h	�Zu#{��Dku����D�~ղ�>��;Kh�7�A'AhF� �l~�-̭"�4u��w䛼�����\�Ò&��A����Ǜ��>=��A���],�U�����,#��xY|0^6��`I}��:(S�}�_o?�i׿g�aO]��@/$YI�:�y�;�/Jq1��nO�`���OA.�ţ�cnC���ׯYע����rs�(���kJ�L��l�5�-���O" H\v:C����O�W�k5� 4Q�R��L4Q$�lJ�ArR=Og.�^K����a� O�~�r�V������m!�j7rRB��]��6=h�B����h)�t��_��WȆ��~����y]�W�@����v�R�Z8�c�vY��H��v3Ao���N�&c��p�?Wa���L�`>���wYu�%� >��B&�7�#a�t����b���GTe��"�z�Ԯ��c�fF���Ӓ堧=dΨ�芫��L�9�W�i7t�9�"��U��M�'*@0g��ݹ��H���(_����.��	!U*)z4g��������#=O$~����O��/( 5{��}�� ���b�}��a5=���+�����v7�	���@"�^Iه��0a����"�+����6��wr�'t=eŒ2o�ڍ��rr��*��l��yZq~'�V��K�����	;�2�.]�5���?���{T�;�UYl%I�v�bu%;�5�m���L��#i���WJ�ь4��:3c��қf�)��G�0]�^�aVT�B���.�J����$�m��� �����L`�	Ĩ]�,w���>�# <��g�4�i�!+���N!��V�q��ݸ*i��3����AxC� �F*j}����f.Ӡ��ZJ��#LZ��ݲ�<SD��d�++
���Z����%c
J�����n~ԁ�|��Z����'���Ţ,H@�u� c���1gkc��%�]ъڇy��@���i���UӸ�r�8�e�(�+���6���݉>�=�:GJ�T�Q ��s��y�%"���K��!�ތ��}o&��[_l �ƞ�{�3ݼ�C�U$�>��^�-w(��j�TG�X�g�k���n�(�GŞ"��=vD���16�����*��f�=�Q����G�F�a��Қ{K���AgT$�B�4,>Ư��ea�:�gּ��7�p�/���`%�FB@�g��ɮ7���k���A�τ�b@XM��- ��
����<q$խ����{��-�KOG�*�x���� "i9?,9��y��H���N����g�^8�D�O�ߡk����~E��	ar0�h4Wa�?��s�vQQ���G���hۦί�~��zp\,x5��yo�E�t��X4w��g����C�"(�U�_M+L� �{t/c�_'7�Vd��nJ�{B �;�^����TN��V��JR��F�#��v=�x=��}�B��h��ף�������1�%��Њ?f|Jq�h2���j��	� ���}_�Y/�N�	�y�g���4#s9y}-B���߭�����u��\�MS�bBδf�J�Z�ޛyL�҃���W�6��ʟ�9�~���;ϭI3��q4�r�[�:�&N�>� �l���Z����',����������%K恠RQ��ʓ��\|�b㵻�d����H�(�Z�� �uB �$x���v��_�Y����^]'��0�v��!�Ջ;��y�T��3}�n�na:�����}�`��ٲ���^�tZ�ΎW*�$ ������OC�J��0a^W�;YJ��̒#��=o�Sy�À�x��ON%��H����n���a2<d��� �m7
�{��-h���Rw�K����e�3���y�������� lfe�n�x*���l>����T�}�w�i%~�\�|p&�jC��c����DE�cL���7ɢn�0��­�a��VL9���{:Ñ���$�λu���v���� O+�VA�~ʳd�B��C����Vo1��j���������Lƭ��ɚ�d�5A�N����o�Z���٥C`_5y��|����ɜ�OЪa��j0·?��aLO(3�Y�@�_o��`�"e�K$���M�L����zuB_��ի��Y6��y7����L�!�
S/���|����M�Ǭ�+&�x�C�:)7�WJH�! �1/��	��_.������FN�@�tJ�1���)Q�\B%���3�V�'��
\I�\z��=9��-	I�z�~UtpL��;���'{D�b�(j߰����Ykغ���yj�p-��|�~�Cm��~��e��hG�0A��Rb��'6��J������=��hw�*˅�a�UyM�%�J�ȫ�N�8LAu.8b�A��[���K�\m��	�}��b����%p�ݻ���Z�~㏜�"�� ���u����k~� ��ᵫ;�r�?5�C�A|=-Me��)���t��)��G�,*�e�*�Z����z���!yb"yG5 �јW�~J0>�"������	@Tc�*%�cl��.̀J�pꋨ����i#�"�꬙=��gq�Ztn�Q�5%U�:gGg|�o��k��i-?��	�*���q�3��_��PX�G�t-��+_���j���N�r�ۭ�#�OʅU�F�6�,<&V{��H�ߑP1@X�%ol����շ|�&L�м����Ho}W�gn���5N������dQU~$ah��dѸI�9Oސ���j���
tn2O�Uc(a�j}�{]⭧�ɷz-���WI��L��c8������)��{�^���,�W�;���1�X͞�k���)�Mw
q�==A��ݭ�؜� ����-^H4Z��t���啫��n��.�""�GW�÷�h^�ɽJ�官�]��@T�I_��B���*��*TXl�9��[��Tt��\��$��$gzF�����u~J� �ϕ�6����.�-�2�65�<x>�>�ׯ�[/߅�A^"�E���2\�vκ�������l�Hr==C'��W���Ò�U9K�E���a���]�:���zi�^�$���y�D&g�������7����%�x������G�8Ҿ��R}E��H\d��4N���A/��R�{T��J>;�|�$�~���F��C�c�`�~,�v�of1K��^���  D�[Kw��C��&���dD��1�k���t�_R����b�p�C��霰��e�T2��ơ����i�2	��- ��� ���K����K�%L΍���!�*H+$V��d25�_�r���h+'H��A6QR/'�������0���Eu����y#���PJq����n!(��"���j��������m"���F��
��++$����	�M*��F��%i��e���o
�3�/��K�����l����a{~�2TT:m�Օ��I����'nA��=7?�����Q�wQ䶶�f��I�	������SU������;lOFi�s��u%S�k����J��:a������,�p���EƊ�����`�s#�����Ëꄐ�~͟�
�P�V-CO�o�o�H��i��A��f;���x��<,��ߑ�mU�Q����b(�h��u�U���c���Ԥ`V�2{� a�T��a�D~ǆpȞd��vI^��d�V�������ٴ*�x2q�IS���x��?N	��p�/i�[u��|���L	����ց8�4a!v㽡�����$�����!u=��5a@��A��v�|qS�;?1�mð@x�A~fA�%�d���%�C$��ȧ�P�=��u�V'	ٌ�ɲ9@�y�u�Z���3M�3�+��D�گG�//���H�z��.�� A�@SB������kTʸ��ч��Y��7�ny胨�$ �]Ѩ]��v�Pc/O���mi0������@R�A�H_f�ۀ!������;n������m��Y��b�נ�y�h�2����6��w�fF,���%��c+��
=�x��*/w�<愈������O�*���$�v=�R�.�����T����ꆼ�{I��ĥ��kՄ�6��R���r��sbdZ�w�����j����Z�L�7:���шw�D4|�~�amk���Q�7�"u;T�7�7�T�Y���զ���U|C�G��8����V2��Bp�|d�&LwL�oڷ��M������R�\�[�-X��Kn1]J^��כW�#���!{V$�p�Tӈ�J�$������{�n5�o%��W[��#*��������2$MS�-�Ld��͂��#P�)�m��ѢI�����˸S;:��{|�Φ'��c>��Z���p��o�T�g�Vݪ�L�E&�$U�M�a�2��$�IQ�k��n��.�����q6^8P��ݫYoY�iVT'�UYZ!��(��Ǟ�z�5��T�"*��5�c��b�^D���==�v�J��ZԷ�~�Jl)D�穐2��P����"|��δ�gf��1�eN%���4�dz���u��@��ybG��N�y�!�ВYL��i��yԉK��G<���\T'qH<cѸ����X�!�L"������/����TUZ#�8�&��#=�Q̯#�^]�Zt~�X4?6�����1��w�W^�hO��>^�X!|��_�$����q#ӄ�������<7�)#����4H� !��y���`2�q�k~���M�hQ4\�҆.�����a;,X�NB�.a��Z�h�+eVl���ܢ珑<�<���L4��7�Og0i(���3_����A���re�ܸ�Hݚ��gUa�*
$ڞk����"�T��uD.ז�޺Z9S!P�WhxV��la�כ ۥB�qR<�oՆQq���O��'H�͢��0��X)���:w��_�NFT�[@���pj=�n7e&FTZG��!c���7�
��=Uc�G\�^�z]
��7To8���+J�2���a$��,����U����,��pB����롡�d��l2�*6��{�U���p�Γ@��2�p4� �����;f��Fe����0=E$P{jzNl|6|~���Д���o��u%���Y��Wh�ZJ�.g����q�L�L�x��[(��.(�0$�隩R?���&7�Q�j�l�kq>��h�#�	U8�����R��b��w��.Xɍ�$�ui�>u�]��5[X��m#��5����8���\`6s&3☪����v#ۻ�HꃟgD�	<���a��ͯ�`rxr�_
6����ލ�B� �v�����O�j���wCaW����W���8��_�1�Z�ċh�PI��v
9!�?=���5$D��gD�2���@�-*��#��{-z�K���bEB)�����P�
E�¯~JXT�D�^�4�O6��ۈI�	L�$��}@�e/:�a�Y�l��tI�K3`i��hRSkk��p�ؐ��KTes�uc Q^��t`NX���~��M���S@�Gc*Q蘾�\�j ���Q����[����9��9��](B\ݮOx���Wӻ8!�4Q�ye���6�S�X��vKI�ǁz��^=fT��h̗J~��-�0���z��k���b��L>���t����y����}����Ӊr���E4�����l��olւR̽����l�2<��k���z����ş��F�}��&뱃��$^ /��U�����^V�Xr\�D! ��}��:#��\T2�v<�l��P!�J��%:ш,v�^	Q[�"g?7`	����-�\6m�*��=�.��Le�'"�!PP���^d�x���ߴ�Ǎ�#���YC(���q	V�@�!�B��yw������q�7J~��&�K;�Wt:��/�]��>V��%w`�n�N���F��Sy]2���u�N[H@�4ҵ+#,}�^�G��G�eS*$�U�r�W4�Ub�-ƷQ��.0�M��(��<�8��/��5���}��**��b�4��������J4����\+I �/
S�췿���^�MZ�9R_�FXL)	�N^�ma��`B�����@�o�%/��נ�0��*/���tq��=��V����+���]s�L<�L�z�Ʈ�Ϫ�"(6�_c�j��B��=U-C�c� D'�i���O���k\�i���gb�>O�|�h��K��8O���$o�/Z���bOHԸ��{_��"�?�I�9�� �1'w��؊HP�ͻ9�c���6���A��Kp��aH(��.u�ttMC9 #i��.0~�?ijO])���e�bZ�r�C�̋"Y������ՔT��Q=�+��F�����'��)�q)+���̸C!�Bѻޘ��NSUJ���bw{�N�٣�����|_��o-���L� #��|��}��s�J�R�B�ܠμ�}F�A�Y&q�Y��L�.��Z��ˈC�D����y��+��9Q����TW�2��d~�'���w�ⶐM��0�@g�Vʼo.�$#��|�ț��>�>�����R|?Ɂ=C �N�e��O�?o����!�|�W�!��)�㴻
z�ٻÆ�^N7�e:3�ڋ��ż�<Gq�"�t��[�km��Du�&��E{��G�-�"��c`��������^;hP� 0�<P�\Pt�_�J`ɏ������aJ�X�~u)6&G@�ș9ѪϏŢ�y=!{e�J�MQ�o`���\2���f�:�wj�|R�Ia����PcPw�{���Lq8�����sb�WE�Q`n�d��<bi���7V_��c^�'Q�&�'b�Ex��#�|䍋�	� 8����n��<c��G��wɘ�B�:����nڍ�`����Kʁ���n�t���b/j=G��W�Qy��\Ѿv|�Ox��b���������Q��,��)����8�DS���Ƞ%bXÐ�qyԆ�y�TR!{�P�G����߄Y��H��-6�w'ң?��R<\�d�qH�u���W����꯻�a[�9/��g��li)H=a�CR���u���y;3�i5��,hLA�z��<<4V�$��|\^���_!���^E�VǷ "u�b+���u��)9 ��'�d V�EJ�^�����S���wY匩qy\�5�C@ ���y~R���EB':QK��E�������%��'� ��ܫNQ����4�k�#�5ȩ�����h���)W�T���mxi��J�JL�RW�)@GyQ���a{:#j�8���g䗞kj�6Ŀ�j�Z��Z���[n��Yu坢OZ��Q9V�k�Jt��.*���x��:F� �,,�C�w ��1ڱ�y�>B�RIM�M�嘯���� WG�O��m&��p�
������(��'r  ��7Xn�B�N˅� ���	��d��V�g#�p�=� ��lF'����#������� �v�9�P���~."~�~ӡ�}�ٟ����25��.c��Mݴg�A�� o��X}�I���;$�3z��
��/�;S|���TηQY]R����(���\�0A����6���
t��k�g}2n��D���`lȜ�y�$��l�H�g	V���w�"E�������^w
�A9�F6ρ\�4�)
�.(�#��2B[)ҷrO~u�}W��L���.8x��
#6�:~;�ӄ	�EUĄ>��Y�'k]�*8�%*��B;ܲ�c3q�"���iΉ%��KS�,�m�����N�/��ڹ��ӿ�@tMTԍ�T���M8�+��n��w��+�V�MOUޤ�~�7�8�ϙe��56�7��xAq�_�jX��չ&�Q��ܧO^��Z���N2�'EY!�?�XBhZ%4qZD�6�o5��ٟ�-p�C'��V猢�Q;�8�.ʺ�3���{cʾ�����]�7;tz���$�>,��ȯq)N�,? !��ߢ������J�j��`�r8��%�1��	ŏwM��N*��]���ХP���+{�$׶ J�������w��]��gG��vd�d�a�Y@�������Q*�s�%�܆N������6�-k�Nuv�^ah�4d��9n=��ϤwK��O���U�\9���k._�a\�Q���Ǿ�DE�_����f<�n��2�-V��D]z���^ڢ�ZN�uO�+�u��A%q'�ͷ}Q�-@Q�}����lR%���U��^Z�o�Ode��\Y�Hڲ�4U^o��?}*\Ԍq��p����r��qJl����}F�2�����/QP�l�֌RBܛ_
t�`�~�E}�՝/-\?5>	-�Vz����m0�M�u�����#�p�P��w�9�{(�� ��_�"FF�	�� |��B��˙2��>Y��J�á6�~
#��	�l�x�l �A,s��k��?��*��A2�?�wf6���nў�0:�-�)y����2Rbч}?�H���Y9$�
|���y�q���Y�.�W]� �F�c*�p��;ƈt��)���U��Be�޽��']�˽*n��J�������O��`H��S-�{
����vD^N�����94|�V����p���r�Y=�~8}��������We���޺��#y/�zF;��ةCt�@)QԘW.*I�bf��ܘ�;�Z.����/���	@Hp[J��Yton�lz�.+p�*w�x1��;1)��	2!Y��x\�9����A����>� n� �F�,9�O6Lu+-��:��󿍪p���������D�Z!��������QI%�ڈ�V<��ŷ+)�탃ǯ��Tx{v="�k��`�:l�A̮�K]=P�-n��٘]�S�x�5��*]���R>{lY�o���]�R��{J6:���q�%��?>�~�AX�*���'UpHi��j��,/�伈�e��K��˝/Rk��4.~��f6Z�.\�z!~�VLa ��=���a.rg���
�b��P.bL��b�h�r���aG�s,rɣ�-�\{��U�3�~4u6���g�la����݋5�x�!J�"KE�x�Q��q�� &}�W�Ю������&GȘ�X��R�t% 2=�\ �{�f(߽XY�Po�S��:2�;I��j��n4�B�SQdo��=���q��w�W��M�^��,1���u�W�9����]�3��O�CԺ]��h�R�i�#�����btݗ��Mr�v�x�'��c�'�,�x
'&Q�e������͎^ϑ�
�c����`�N�D���E�Y�>I�j�N�1{����`L;۞,��t �׿��p�=|m�T�3gd0�Vu�(�R���6
cI*v�2O�Ukl�pV���Z�1q��Mw��i��-W��M�MD���o��~��#����)�rb<k;�|�g����8^�����r�>_ >�L��c�S�m����Au�
��z����~r���\i4P!�s�->O����M��]�����r�_-�.)m'5 �|Y�j���.I)�hy�v�}�;
ƀ�R�:��C���7��Z��YU�;[�޺cC��*M�����L�e`\7SXǯ���2�s��g��f^L�Ѫ@T�~������i��s��[�J�!ESxqڏ��x�qe�_���6S���O@@+�F�uZ>���)ۏ~.��� ���'��@;��Z���<����1���h��e�|����i$�{��>���W�G{l"v�@<�WŢ�8�{��~I��$�;����e'c�/���&4�(�!?$�?�͚^5��܅��F9y+���={Sf|7ٕ_��g1�a��	.��D�6��ㇺg���kzf'||~�5VFvx�(��*j�����5wH
�\%��Ŭ�eMm��ݽ?�V#I��_�� �|U]�%�{�VxH�<Z���������<)Gx;��zm��w���>�=*��Q��h��X�*�����!a�Y��U�=�?T=�{io��lٔ9����q�����}�!�2W�ΤB���0pj)��!�&ya�reb������$�&������"�3h[���8��ʚ�����ڒ�s�VW	Z��>�/�P�$�sf��{���?&��P=��r9�ϡ����Q���E��e���dŵ�����x_ݳ9V����tH Ɇ��u��k}sc�3��'Z��Be+��+�.��~�Y2�L���	���G������:��%X���ݕ�5�;s�2��� B�]ɯZ��`�{$͇���:#�����~%�KOIO50֐x��OBwh�h/QG�΂O���>7��cF�&����v����%�t�>lQ���N����?_�E���XŸi�B^��I��{U�9����5�Y|��x����o�Q%��<�''��&vIMl���9��>3�e	ŉ��LN�{���g��o�(�\n�7�TJ��ltM�R�K^AWӟ�h�N~T�j���2�X	��"��v?fv	��\/�9�7	(�ߦ���r�}�/��f>��5W7��.+A'��N$� ��I����yӾ��K��9��ӦT��R��߳�Rތpw��\���8��1早�Άk�<� �;#O��]Hh�Ţ7�1���K��J������ ��FJm�u��w8���RS2�%���X�&~��2((Ϋ�=�+;�2�	�F�x�xjK��D��K4y�H���O<tK�'Ip�X��f��Ϟ��>� ����'����,��el兘��j��2�C���)X�o�=���m����R�R��Lҭ�*����!�iL �)�}3K��B#�F�6�B;\���3�.�M9���a��*1���dY�)d�{R_����*�P�|1�L��e>GO����'�`����a��A�����x��p�[Z�򲰰��i,1��f�Q�RJ�{��1u�袑��o�w�S2�ıl�O���zO�������V�7�Z�VZ�vC.!�ڍ6���k�.(�H��ڸr�^&�Km'@0�T?;�?��_ٷ� �2��7{�[}+�1�N_]�j�v�P���;2����6�x�9-�r�a�A:�W�2n�=#��W�����|vYvğ� ڻ�Dz�e���pQ�-�R%pEE@-I1"tƊ��6ЕR@�Aݤ��O�;Z\m��@��`�j�y��s�Xl��%�+Ŗ���yx�c`�c���3�e"c
u���ڡ��<2��x_- ��(�+� ���ӱkx�V��,��!ϩ�]�6�Cp��>̴��sm��>]�ם��3�@��b��j�mY�)!��ǇqCQi�KMd�M@X5���Aqߍl��Q�&�=�(�;|�I�5��|X9��؃u0�*vB���D ��J��!RU5Tuph������=O�ef�g1�O��g��|����v��{l����t�s:��� �y���ds���0�D�'���/_G�u>����·Zz2c�|��m�9��"��r���Y��>�y�����n����N�B�J��9�L��NҚ�̊�/�G](��m��4-,�v��׵oS������|ܑ!�:C�qs�Pw+l��/���r
G
it�����u4�Zq�TaG˴C�-o� ?J���Q@~H��U�����b�
0
��z��k^�18 H��g�O��X�:dy�^�颞Y��j/�ٶ�/�GI$cຕ��� r��]A��8�C�(��ș�\X45����amQƧ����]��".�R�4������b�X�}p'�\�f�1���t$�R-���'r���;�%�����Y�.p��֍�d$�G}� :
�Y����s9�z�������6��z�w�����_����3�. @�l���A�իN�[^���9���p�
t2�y��Ӷ�{�����h���&�>]>����5%��೑�:M�C�C����O��z�2��L/�eG�>�c�x�U�ό�d�ՙ���\B�ǔ����!�	M$2�/��3f���H&�ӄ�x�B�TL۰�L���,t�ϸ�7�^5�Q��/z.#?e\USQz��F�Vзd�+�PQ[��䫢���c}�BY&%~��b�&o(q�ծ�T�-S�Ac��=��^+)r����Wu�J"�Z�n�� l��8.��z��"��S��@�k��	��=��c#��ݭ�3�U����h����s�d���=��w�O�Cڭ:2/+��0��*�^Ճ*�0�Yz��ጬ`.o����C�Q
~֜�3k�F��<��I�r�LӵQ �s��Z��rv�B��du�W�g�K�i}�������y�����sg���z��-�To]���_�=|(�=4揱MX��	�w��h���;ϙ-���;�%�6��k�"�K�����?��������qU`V��S����Ct���B$guK
S@o�h��z"����B�ĺ��*g*�^�M4lTҬUtGē�8�ɻ��>�C0A�W=(Zo-3�G��/k����,�H����5�����L��ޢ|�͛d��<o��H�փ��ٶ�ί�sڎjD�vI4�󄝕���|��4`�y����Z�9�d���$�B޴�Ч]{���hâ�WP4�	{�/^��O�B�x�����{�G�(�K�9�uP���AT��I�h{��G�A�W�%j�E��j�IN#�ì��.IN�4�D5*��h>O|��	xP�pne�(�9��YU�w�J@����xxY��ϐ�4Q�둄���&{�jhK�
��	<�S��?
����$��C���h�k~�[@��'ȟ�u��YQ���~���#m1g�6����ޱ�9��B�QPo����T0s��wOQv.&�d���ǂ�!as>o�<��c��Z@���t/������Q���%��?/K���uſ���~��]I��*tڵ��^_�(��hXD��(�h=���i��b��M�9��8�6_2�u�S����t���.�'�I�cM��9C��ں�/��ǭbfRm�|*Փ��~��yF�z)[���������t�Zz�Đئ%�֏������:���C��׏�8J�32r��H2�r�}��V0���ޘܣ��Iq�#�3&nYX�Lv��I��D�z���rh�����-R��I;M���
���I� �dM�
��V*1�������sas�
��(��S�eCݔe�/D�����P���{�d*�7���X�c��ˮ�3k�l��1�~��M'4��C�V4�Ϡʊ��m�l/�0Y�Y�}�Q2����^�I�y�*C/z7�����b�,n���.��=�J,�c��D����~9�j�������X��Ɉ��m<�7��}6��*��a�*x��S
:��z�y�g�K���C��G��۝i��\�Yb�>=w�j˦~>_����i0V�p�'?�!�MJ�`��[W<�K�I!rp�
X��\	��Gڟ<+�>jNQe�����*�C��]6D�G[���M2Վhu���K����0� �U�C�M?���3�t@E{��Ȥۥ��k��U+{��NYS�3�#Y������bu��d�d���o<g�®w}�����o���Xx�3���0��X�4U�a�HdF]�i��1q�QL/�V���1�$3��an���O6d��n�!��:_��$]�uܝs���� �#�o���H��{D�)��5��ޏ��p*�]ck��J�)�����[(�{t��T�:�|Y����B��D�9�d�q0�gs��S8��PR��F�u��ĺ�Yb(�~�/����9��R$�Q".��j��ܟ�BdЈ�%j,�\aյ�u֗LkH&	�o�n���x Y����*eq�}�e�[B�\ř�����WIq9�#\�Ĕ������+<���g6�{Xrp���&&J���N�����j۹
=!y9��-�x��>���8�mǫ=Б�^2G�jY(N�>�C��D#��7|UM���@6�[`���y���Mf���?�l�J�Q��L��y��-���P�7�w)�B���|
	�Q&k���x����Vm�#U\.vV��g���>I�&DD�-WO���.��Nܗx�eѸ��	/���R��,[�p�B�~'��0��;���鲺'>'0nk���xA4#���+���[���2H��5qֵ\�u+����^�:qw�߾�V�2���c^�C��eYː��C�֬��ys՘�|U��ߊsM�-��{��x�� o�P��@Ha���m�T�WM�̫�}����_{�(2`f��C@R	 ʊ��e*��xC��x��Y��O>�I�[�Fm��XB��@K� 
@Es]�D���x!�I} *�i%���`y�κ�R7�ΓIK��ٟ��cA�ՑVP���[\k�y�$Ӊڝ��T��������K��(!��J�X�W]<���U��׭��#���\޳y �����^��(�\ru�@V)[:C�Ak�9ËF��/���5QF�/i�ׯ_���k��X]T�Z�4��t�	N�����2�yc�-����j�Ⱥ� b���y��Jn�a��@���m�}�-��c���4Z����BGsK|"E��p@�rV@~�1�rpF�KE�z���ʰ8��]A,�� ��-�Npww_�$�$��w��]����l�s�_�y��_�3����Uo��]�N�sY���8�0EF����@m|?n�/I�v�� V�H-w�ww/��9���2���8lI��=f��=�ۡ����J(��FTei�N!�	ˣ��~.7�)�T�<rGR_[��#Y�U�.Ȱ��D�ey<5J��X�\�3:c�0���D�1�A�8��
����c���z�Ӻ�"��v�sJX�/�8�,�[���Py!;�/��Φn�o
fB@�"9_�M�P:Z���6��]N�hT���}oB*<���/� +��Z�~��g��}f�m/tx<�����%���~)ph)����F(�Y��+>2��Fލ��I�˜��^G�f;�ȴ����U	Jځ���am5��^��y8��,j�������M��X�y�5.��piQP�V���:w^�VH�G~�Z�K+�?������GCjض_�=ޖ���}�0n����
��fU�ׁ�B���Q���S�c|�$��Y.���*�3/{;m�E��\h����n��Sz��SCI7.�2���<\.(�w� ��>�r�R?��=i�
�=�UA�:*��j��D|SOGد��=��T_�bXCâ�.Y�P_dz��<�'����y�',�|{S��G �l2>iޛ�(~�h@>ܛw�q`�j�n~�Ab������h�iW�5|��;`V�k���!L�O�̽܌��W�|ݤY�)(�P�~�7Mv�/&/5�ÕY�]K������dL��rSR��n�>��pL+'�lT�c2�}C%�gk	���H��2�6 �var+
���!��]5ɗ����/=���$]�3�����~#���t5
T�2��6����H�6�V0���P�H�C�Jb_����;;�!�t�;��4cb�`�NI�rW���E���BFbN�X��K��}������U����~�{&ؿW=��
e���&<!z�(��S"��}�z�<��M�l{Wik����u�>^�4�֧�Y!��9ޒ�_µ��������e�Z�Ǳ�o��b��)~am��"s�7�����ݿ��W"���NK&�V��<}�L���0�5=���G��+�b`0�&}���i�χ�/,��S^Cᨪ/GiT�CdJ��~������d"S�r�yj�Y@���6�r|t��S�lV�{k>��S�+F��(��sOVI��:��.`;������_E�DM�k��E���\_ļ㐕.&�,g{a�bN%�񧒥Q��П�6�١Rr�F�渤b�N0��� u���L[1h>P�,�%x/UЦ?��X�;��@a�h=6�VQ�f�֒��&��3��]��Y��w�y����KeJ{z�z"˧����!62�3��<�� ��!/���O�rf}#¿�ƒع����Vu��KV����v���{q%{���WG���|]�5���(*��q�J�>[��-l�)g:�%^���"�$l��\(u+-�k��fw�1<�D�P������6�݅2��y�ļZ?q��ե�gX�S�H� ��Km��������Ŭ�9-[� q�q^V~�(қ��D'�&S�,ۊ�RX�B��K����<Y��`���1��m�)i6B��#C�Aw"���B(�bg
�	-z�h/}���?�W�Xq3�uOq��y�a��f�qc4v�Х�Z�5d�_�_��?X�������+��C;i�<���7��J9��?#���/׈��܊-��E������W18�+��l�o� ꔃ����]�pI��Q�}A�t�g�"k<D?�/�.ΙP�c��QT��:
��MLf����W;l�-frl��?rbȤs�Eֲ'x�'���
������
���X5o�ךt/�y8'��!���fh0��a���݋Z��}�¾�L鷨��D.%��.A�%%,1���N����o±.���,���1�6fo��+��^F<��L�(JEˑ?��k_�
Tv�
��{O�)����_�PSgG�I	�$8LR��O�Jq/קaO�/���/BL�ͨ	��7���PM�h:�U$_C/��yC᧵��ח���Ӆ��&��@ ٌ�����L+�����X��3�Gl�Ʌ+mL�X�&�����A�2
�A��sl/��;V:�`�Y�X��W�D�@��o�H�V��/�V*V*��X���/��g��"2���S����aI�?+��[���e�pWj��e��E̺x��p��*�>���*K�ϙl�B�,|���
:�7~SA&�p�8��g�jX^��7��|��Cb_���c�|3�O{�oȤ5�i��#)�x��wL&8a��7���f��F��,*9�]�p>��3��i���u>vH����̋��4��	Z��/h,1΀�eE�=<�iִy��t����)�k
	�E�SG���^�Հ��@}Z�(B)�xn�����o��Pʟ�:�s�Z
�ń�\�J!����O�4�PlmP��ݠp��-d��'��v��w=u]oC(r�E�:K�z嬌$�'�[�2��ٱ��n~�;��T�,�� �*,^h��#�qȆ~j�G�31��n��+D����Ӈ�T)���Ԏ�^��S���*��.��2.�j8�.��j�<�7~�
�(+���cU�U�0�cӊ�\1�rµD�/����U)�2|1��3B@299٦	�}�W�y[S@斠KLMK�� X�=����n���K����X��IV���4U�WABٴ�>�ȼ?��a�'^�O_u��&�k�qfF�"pMyT_���>���`�5k�45����m���\��_L7ov����2�TtpW[��-vUw�w�3>J���*i�_�� �QWK4Z64',��I���=��g@�	�J4=X��	I1M&8<�)g���Z���/9��Z�)c��u2�ӵ"g�۰F�T.%�%���*)�?��)�<����3�$���3,��iE�[ԧ���Y?L|�'z��/5�i�����:�����Z`��YjA:,�\����FL�cZ�\J�$k�a3�g���0����k�!&�x�Y��j]�A�9��-��H?�(��NV�a�>F��#��nԔKIC���d�t�>�����c(a��o6W�Sx��=�3I-�,i���@֑{2Ij�t��`�{�5v�1�{͓t��j��p��������)�(	�y��4��J��r��9fm�Eb�B3�K�C��o#�D�X;O���NM{Y���6:�
H���~�e樈�0� <��k�Enm8�Y�UXO�@�K���k�&���(��[���l2�ݩT|�V$s07�B�3j$E3����V��D�z��2�&X��"/�x��¬3�]�u���/F�!�ۘW�&�A�I�>�gn.<�?G�,]��URr����܋zR����:��&E]G��b�ݻ��F� �4��%\��L-☧��*��^Q��	�0@j�~�7u*a�k8�L��'�XB��(�
|UJ;�Opt6��u/-D��NpR;�	�`®i��2\�F�V���/�H����oᤍ��Hc�y[�t�U8�"���.E�E�/�K$�{w��b�e�a����������ʑy�s�]��Q�r
W	Y���8�������d��_d
#�k^���+��Ͽ�KiLw�"4>�ڛDp.r�� 9m�t	Y�PzM�\L�;���=�45�0���rz�9��|��Fv�	LA,�~�<���qo$�������B��A_}�^�6́�����d:�+��~��ɯU4�Ue%Y{�ks����=N�N��:��/o�<�x̸DS���~�=ɛ��>�1�O?�[��*��"Q�5�P�LgW�Ǔ@��+Օ��f�X�w��
�b�#wC�X���"�C�no'0�Ԫ��#����}�P��_ ��4n���	]��sK2�wFF�撽�b���^^�۸*��?��ɴ�33�𺦤� �m��?������r0�$��Wg�E�wZ..�&���ܯ=�3�J�t�o�*�n|��D=r���A��p؊\g�m|�3ݛ�0�j��xO8V�I��Q� ���[L�������/Glձk����8u��&��k��بcH��h��*H<��Ez��oU*���l�
�+]�I�x#�`�
vK���A��)]�e��63��<���v
o����+*W�^?X��ð�����c�qU6U�|�n!�@h;�P�����}3٭:���<��>���Tw4_�����=�'&`u�g�Z!Y�w��h�&�J��_����-\X����{������`6�BHREQvd�܋.#n��hb��9x*�p�,,fأ_n���;�\�{qL�U�'|��ůA4�ޜ{΅��($3��@�b����[7�yߙ�x6u�gȇ���J@��'M�=K�T��b��}.8��L6xϭ��d�����(�Ԡ����4d�eF\�=eJcdPE^�y��;����c'�l�q��SF��apC��W=�^����Ļ �v:�\�7 q��ɬ!���
A	�r)-��א��$d~���5ء^]�	<�Կ����5��W�Ԝ�?����[pR�AN�o�WR��U������!bz��؞�J�0��-��
2Y�o�u�ڍ���2%��jn�,͢N'�С��8�e�|1�7#qݽ[�[ցE�3z�1�r��Ig����Nз�����I���+��pI�7\�zDڸm?�f�R����>�N��A��׋)ԴBT֠��+5�r=j���u99� �m&_j������ľDĪUi`�s�֣�}��@�O|F������M�Z}���F��F�n^����~R�fE��.b�qI��ؤ��z�:�_� Ib`���ʖ^�V@:�m8q{�X��� ��/��be�KH���T����?;��E�ލ&���̣B����]�w�2�T(Ϋ��g��Ϊњ4�͟��s� �����{q�;�o�����\���(Ń�D��nB1��h���3n�뺘��k�<�!5�>�ф�+��~U���T�x��D�g���I��Ƒ�je;�\����G�u݆裳h�[�U��	箲f1f}\Bk��~�t9uɲ}�c�P&�����*���Q�O;�ouaEO@u'Xl�L ��ȹ�:��$�@SHՏn�������J�w�$5#��T(� RYK-8�@�F)��3�zN����U�%��$i�<>J�ˮ~e(w�[���t_�]�i�-E������n��CC�8�5\;?��bw͖�Ɗ�b��yݡ[ ���[n����L�Z�0!2�k2��*
d�+��1��O��z��}�O�2���`��T���#��]� $5�_����/�X+T��t5m��ȃ���t[4	�����A��-*���.�m�?�s��o=�.�o �ڔヤs��d���v:���-��پ�[Ӕ�v�b�FY-����uP�qn�.�3��/@.����",���Ϟ�!��2�bUW:�$:����/��T5P\^(n���jN!�cs���=��ԐʲO��A������1o�V;�'�>ŏ|Uے���F�V����TC��0����f/@X1�X�E��`ZyIě�m��F�c��i�9��!(��oZ���_�8*Z���ň��Y��
jTG؁)h��o֛�%�E+j�ͣ���d\�n'���.d�N���?o��Ԫ�?��I��:A�B��#$t@{;	�B��!���o���b"2vG	;nVC�V��1�d}H�8D��>n1B9�?{��>s퐢��h�9曈�k�zn�~4֗��~>���pS�f�Ppf��_mG�}���|��2�?�ٛ�9b�H<[,f�I�)#wT��t�<�%�ZH�r�=��� �������+�`E�O��T�����nB4c���O��`5Ą|���I�J�PR�%e<^q��џD#���QKg��K���)^WBQ�pL�z}��vD���h/��� +	��UuTw��D&�zs �R֦zVG�a�ߠ�������3%�5� �Nr��=��`ыl�&��C@ؒ,.�b3N,��V`�3ܴ�P�W�H9���ʗ�bfN̹�m����zd���	Jh��X:��9��ǡWƬc
s�w�_���+������3x�k�^������i���+ap�,�O�Ե��9�tiiv�x��M;:���7��"�˳����6MM�4�y��v�9j�μeX�ğ�087k��*���M��L���4�/��c��f_�����<�R��!��t�~���i��qG\��7wa8]<�P��#�BY1"��/!��/��CD]O\���>Ű
�6b�1�R1)��*s�p��������H�f��y�I�ZJz�X�`풗Z�#Ò1a?�1��]*�A���s@��8��Y�h}�O�ū�z�	�T�F&��!D�4-Pߗɮ�O\Q@��A�����E�G�/�6�=|ņ$>g����McD�����~ݨ�N�� �w���<ܰ�r@�x���Z���V�n�.��f��Lp���$��u�}�펧������r��ܿ;�(����l����#0b��3�<��-�"��z�����(�b
�����?���ܼ��<��^��f�%Z��BU (Qٸ���|RL(��"�J�����\'IOu���>ֻ���HT@����]������g�F�(#�t�Uq�.z�b��|�����K'���*Q�qAD\�'S ��"�ʅ�XIT?~D�R���۠9Kbʋ�j�c�!E���ɴS(!�@<3ؔ�������-�7$J(o�2��y�ff���?����X\\$x�@\F��B��;�;�ݶ|��?-�s�^��n�����"�������/gLy�kE�۪ݵW�no�[�1Ƽq��?�o���{��=�6\f=;����IAkh�\+�6�rӎkr��b�S���m-����-6�Y�o�i}ۍ����|���^n]�EE�|��?c>�������H��t�oޝ�Ҙ;�c~"��9������#���JI�����>�����Z����W���T��;,>�t!�2��%{=�H��Y��<׈y���#'�)I�O'�x�_��0�.�N����c{�
��6J�ޅ���:1�p��8~\O�����	pC�Q2��}�|����q�����i����w��߮8��ӂ��w�jʂ���*ug�S�=��\�G���iu{���l�3�e��������	0����J�f����ӽ����<�U_�kul�K���mŖ>�jp�pC��H�Ւ!��M�ݏԑ�/	3j@RR��YÌO��C��k-;S;���@KZc���\��?�������gF���3�2��.l.K����Ϻ�fl�ש�l�~;�]lmŵ]�H9��T74|ʹ��%�<�Y�J2-/'�\��d��Һ~�]R�4�~��&7r?��N�q�'XjP�rԴ^n���2�����.���a��<�>����K����N /�����H�|�f���nO�	{r�Yl2�|�]o���+B�=n�4v���Z�bf,�[����H��[5�Mm|*R�$]XrL�J��L����3��x3w���<�rki�Xs\o� �>�xwQ���o2��Z{ᖊ��xm}-�|q)BbY)8����Y$}ﯝ"6�0�O�f38�q5+�J������`�g#+��h/c��?#�>CO-�hz�����.�Ѝ~f���.=����Ip���f8g�0�CU��c��T4�N��F�Gr)c��A��g��RҞ;�%/E������^�<�2o��_G�<gt���2���#��rj/�ۤ����՟���bc|G�B9~z�d��sr���@A��i)%q�k������GiI�n�nv/|��	]j98dw��*�ՄE���r3ׁ���K�y���ʑ}�!:�;a��Y�LQL����:�|F��>�^�Ї~����|�K��f���?���mm-꼻OR��mT�Kh�q������i��Y�!�=o�[�}�jZ�Za������k��^��/t&�x���H�ЬeX�2̚�;zH���Vv$!� ϻCr5�J����\"�H�f<��?�nClp#����*Ŀ{^���O��=ao)���/�7���z��UDg�����l�!=�ӽ'�U���&+aE�UH�D,���fq��l��|T�C��6*�ջ֕�U=��<	���O��Z�pEqQv
�E��������z�0����J<�m��ǃ��E�}tt��>m��1=)T��z��C]C�����&S��rŝS���`����l�q�+�@=H��UҬ:2�j!e��´��X{�{V����\�>����h�� �>f���
���\z�Z ��_Zi=�|��#�MH����\\?cc�5��5oz~�g��Q��R�!A�刌4o���֘��]�➞���+V��F/&iҦ�)d׎'���nNaNQ�g�VI ���8?7�ݪ	�	ڄFzz2-����Gz����c���R���9�gzx���7��]���[�=r��G�
�i��PIj�z:�#qe5�_���k֏"�f`JR�f�9��X�%��֩\=�-�����3!'mS�u�:7;40��򑂉�v�4u�iu���d�t'\�D���ޕ�;��z�\�k��{Ȳ�������X��x�ՒHK���3VAsm�ңr�٨wխ�q�gd�?Q_��ˢk��eZa������f@k-�p�^��ƆG�ڇ,���;c>ղ��Xx8�'��2M�?������ї��\�����$Z��<�x8@�L�U���ɒ�nObp�Wl��r����G\yg�m��+!���'c�h�~C�����Nl�����D�u��D��Qj%G�f&5<��ƤB�=S���w#�ʊ�+��%����p��x�������y�ǩ��?m�`|
\ȢM ��g�mu�<�FFɊ眫R�������x-�E�@c��cH���S��g�D5�ٽV�w�Iݒ�"��o�{�	ϗz*M���f䒆�Ӕ"����vzAO1�dZ��Ӷݰ�@�/_�N|-q�N;Lup�j�� X5b\�?z���F��0\\S����8�v/�����6��P�A��K É-�E�"�0Ć���p�}���^)�?��mi�LPY�s��S�Q���|�Xeme|�6� U/5��e�")5�o�����8�ǰB����V�[V��3Z���r]`���E��X����wN=,�h���2��Ο�0U6����R�+!�%m��&T����#3���QذQ��wNI�Ab�l���YQ�>�w�9�v��Ig�)Lsͅ�7�ذ��%wtR����s:q����L%'��^�6g���w��1r��1�X\$�MW7A�z>X(�ͤ:D���ʽ�=L�!�!���C�S_,����Q'*e`D����(�\�n���c	��I������U���x
-�Tٷ����P$_a�%lȧ������\=$���XԒ� �Z|�6�,��D�4�/�~��K����(��x:ѿ�?Ⱦ~�1X��n��ؙ��0\`k8�cr���{C��&ZZ����,|#�C�4;���G�v�fq�s�U ��W�{>��O�ҍ��[jk{q��P����I���@����!(��A��{+)l�5� ��m@/���Q���}��y�|��J!'�7z^Y��
I7l�Xr�-A==b�I����*�\ډ�5��sΩ���2[_&�+t2e.�h.�$�t��^x,+�.`_��(��YiQ�S�+���{��Sw۩{�nr�����S|
W��?�h�=u�ٙ���:e���@���e&de�:_���3��B���g��Z�1�V|�G?=�~��t������c":/�������X���h�	t\Ur]�������%E�f<l�*Y�\�2k����{��$@�:�����1�7���F��..��虏�����0!� 1��y�a՘W��xk�m��q.�f���r���lOۙ�0��5髄�O�,�&RvBTT�d�&w�̙���B�E��-P��8�M��6L��鸊�|����"b����4.�}`f�~��o黊������V���Q{����)p����A�=̺�Z�����=y{��}r�H�X�8dS/�N3/�zZ��t��1?��x>ί.f�͕ǆ!�3���5�6�PCD`�������U���Iհ�W��~�A�l�����K�~0��cƗ;Pń}�f��o�8Q�+΍��UهjCLy��C!+J+]�Lq������E��������i� V'6SO\��"�g��1LsæI#u;�}����DQ�	ŅM=��-�԰���H�	2� S�o�a�d�h��i��c.��J��,��&w'��Ҫ�W|﫺����t�����K����8�c\�+�Ӑ��Ì#J�[%�l�6�9.�G� ��Y7�C~��>V�_"n�_'4u,������'���1/���g3]1�=2tm��k�B�¼���9%��y|nc��_H����0�����$���� ��*M�!&:���=��`ix�l��p-&�����K,�2����9�ذk�f��o�����Sڂ���a����I�n[aV��k��t�X<`��Ielooα�4��a�_^��D�0+�+2؉vzk0�Q\��Z6����
��'.����T
K��@\�w �&�6�ĳ�.�at��,4���>�/�-�bκUMz��W��譡���ht�o���Q��߂S����lg�N��i8+8�H�e�]_�b�J�#Ut����'�ʪ���=��������*g柜`�A��@׏M��amN�o)����q�:��P�Ia����b��w�9�=%l���2���	*���|_�a�׻�R�^��]��}UL����Ꟈ��	���iq2�� ���sY_*����K���E��wwd�"N�}�.zu�AN��UX- ���R]��q�a��s�U����}�0Vh(S|#�%���RS~��/�&j��������k���q7\���6z���=�8�a%� �*�V��+�!�m����<gj����9]�Dj��'T��ߚ?���U�g˽Ȇ����O��/��K����x)?/m������[��l�&n�O5�~���r���a"N�AT��$ĕ��B�EW<�V>��`h���@��y�
{��Z��!/�>Nr�\d/#���~[<�Z-�,!��R>�2@��,�������4�>%l����|_wv+%eF��	(�ae��iݰq �9e���,��M+)sd���,��Sύ���#�{��
��E�C�ݯ�k@"�� jpaOdGi2d5���W�%���j����)� ?/���G�O&X��j�1��HU�P̪pb�!H@^�t��Y��mA��m�IBQ�p�������?id���CI	�}	��+[��"���h���r�>B�$4\(�٧���������.�xD���6�z�u�� *���,b���ё�W�X�;u�W(V�u���g�)m�J��`�aƝ����^^G�k+�+�ك閵�*vFXG�J.�))'��	�'���p��E�W�)���?��@$� ž|ge�J�
�$wlW�d��*!	A:�䘶''%���c�A:�9(+���m��VsL_��A�bډh��? ˰�p`$M�����Գ'=@�b�r]�J���8d�P�t$DZ#�J#ɠ���J�羱��םg�I���0�f�{����=�á�}[�/R<����)''��n9KZ�?�H/ 	��M��6,�=�����Z��~��|^h�-�\��tw�v�4}'�dø�|?�]�H���Q�i�H��Ks�%n�~��螼��B�&�+��ǘ�oȝk�"���	�ސ�J� �2��m'���pO�y��n|jX���`��?R����������m�g�w����]��8���Z��N+��#�R;ܳ���0f^�M��;үԎK�� ��\IhJ9>��|$�x��7t{Xɚt`|��8̦��+���%�ve�A�gJ;
����J�צ�;�T=XK��CTu�?�pH��{�*�b^�y���������b@�8�J tw�ɥ�.aRL�D~y��h�'�Z�)��aj\"���Au�i��K�Be��Z��C��?��v����H�
jx�[%|?�G���p�ni X��Z�`���@�K�m*�f�Xuq&8�+����d�%���3$��<��`���QO����kip�b��TF՛�u�Iۯ$59#sJ��]#��X�;����Jѿ��0i�y@K��H�Z���N)�:W���_6e�©`��K���b�}������Q���.t������F�Ti�]��i���R�l5����~z�R�VX�mde�M��<7���=�V�*���w+��:8���x�X3�Y����65��[��b h�&�"���"N���7M��@r,f�J��n;��9O�n����+�w�d�zےLvÿ�aѐ�H$�n��e�/wU����E�:��<W�p:׹Bo������Q��O1a8L�ηA{w~����mKu� А;q$��##x�'�D�5-��E-V[_�(��q;V"'r�CĮ��jg����>�fj��Oy�L�?���D��3��!�}[c�5s)�Џ�jf�t]�lΊ��O�L�]�?�`	s�q(�����s`���k]�*���d�����u�ʆ��O6O��l�*x~�mzg5�"I��|�$�+��$
�Mq����������p�|[���{��Ipi�`;���(�V��s-�������I�s��3�����b�ڽt�h	��ޤ�oNaA]���R���
g
���8�*�����	���,�w�7E�b��r�ž���_+[�q�lѸR���jZ���n�@��K���s���+4pa��}}�U����^����v8v���Lk��V�/+�$Q!f� PK   Ʋ�Xld^M    /   images/8a38ea7c-aa1a-4e70-97e2-d2d1d9cbf557.png�Y8����Ν0�)��^i"
)��l3�M;�D��Jj��e��֖Vo�C�ݱ}'�I�t77�i�mS)�(�&�q�y�a���v��>�:��<�s�����i��%��F�����B!��dE�J���%�ϸ�|�Y�&�%M��cº.X�yEe>�7;��=1��U�O��4_�q�_C
tLk��2c�Od��|�0���o�������E���&�N�l����L�v��KY��"ڒ�v�9��u)r�W�D|��۴7A�\�kN��pv���H�v�N9^SGK��ӂ��0�i̢S�Yӄ���+��Q>b�?�7��0ajz�!NS���c��h}p�q��e<�Ǫ�Q���\�r��u�x!^�� ʉ�^�]^Zl�0s�U������ J*�:�R�|�W���)ף�����N�f�C�se��ˎTC���Ro�s���	+˖S��CI�_L4w�d�ׯ�荸����2�,Z�y���#��Q�J=��O������8�J�IRc˫�(���~]O���u���d��������Um���K�y&;wE "�Ncbf���X�m7wh3����V�nE���H�� c1QGޯ�q)�g9n����}�Dh���9�����5%$��A�hZ-z,=vْ���YLCD_�U��/�kJH����>�I�f¡����MSCN����)���\�EMyk����_qM	0�i�m(	�;���_Wc,�n:�:�ņK,��t�r�[����
��æ�ݠ��`�s��_�4�8��c�6���o����[�����-ko2�suc�j��b�RQΖ�b�sjƖ� X��|��<L��-AM��rj	 s�� ����r�be���)<�?�I�a(n�܂�ג���^*3e�������䇗�i�	�,)�n�]�r��f�m����ԞA(�%�� ��K�~��
� 8�� z��x*�)Z�B����cqߠ�XD�l4u,�� #�Y8�3������qX^V1�l�r��b����[T��z��v�i�<��~�}�*}(�;�ʬ�/��Ѷ8S�cf��GyJg��i�ע�~;=�"�����;�j{�uHG�cW^�H��s��-V�i�o��b���S��D|mm�%�	�Dt�����V��.�O@{��&���f�]�T"q��J�o��� ��8�A��flG8�Ȑ.R��}�� {�[�5��7����'�31a�$ �	�!��X��� �<J�<m�W��D��W��LѤ!�����A�x���������=�a��uW���h��4"���(��$Rx@��o�n1��Չ^��uYY��6����`��^K ��!ɮEG?z')!]��`/�t�a�^�6b"}z���� ���_��8���I(gme�v9w�6 F�Q8]ӊ��f���@�}�VP�,ϡW;5���S�T~�ߛ���v7 ,K�D^�D�',�E�y^f����N��KlV����Z���Uj���N�j�����$�ߠe��%|�����y��*�1eLB�U/榝�a`�	�� #����2ŷ'�ߙ!Ot� {d	W��� ��L���.@�e<�S1��Ό���� ,�A\�8�<�%��b�%�����*��;*��`��k�B�*
��d�dq��ʈ<�����.��}A��5��d��s�yx^l�B�r�
� Ҏ���0CVM�Ȼ���?3���%�<!�F��^U�+��j�����uߙ�މs�g�g�C�X����]���R96Z�ؔ�W7�rC�7?�L�`�St���[=���BOK)�]�!� 0��IR���rg��n�d� M�I�o��:@O����o(��b-��#)]�/����/��/;�Bqgg�L�5�Mf����Dt�_��WOQ��T�C�3���],���JW�Ml�i�1��5��6HH9��u�w[�: ���UE���a�0��-��c��#�Q���-#+�0i�G��{'���l.��F��J{���Z��)KZ�����A
�w��h�ѤU%XLW��l��@,�4�p�S�q�T���_��P��pG4�شn��q�{�:݊�-��&������F'VHBH�4_|�Z�,g0J(�B.L�3�Lf��<�zj�|��M^=�/k+6����m��L��Rb~ݢ�"�ek��&ÑJ�cXAQ�o�P �<���ZB=������,z�(mRrj	7�������3!O����Pײo:�1�Qy�Eq��`ʼ���Mb��0ϝ/���`!ԧ#o4�C�v,�� ��zU�z�����
6Q�?��ܩ�#d^�(�K��D9��y#^��=��QhTV�����O�o��J��L�0�M �iDy�Z-�w�ݑ6�����m�[_l?�A����k�t��7�lMy7�rtli;���bw�|�?P��F]�#nrQ�%�j�,�C6<�1�ͮ.%��2����5�2��87�C����n+'�)m�Œ$�f��z��`bH��ƥ��2�����^~����(�fz&e\���Ep2��{����}h��h�z֢�i<�U�#�V7A�4�YO�p�OXeb[4ǜ}�����?(*����K�����i@X�*��{���t�s�t��bش�6�g��
\]I�@��C���N�_PZ�D�s����	M��X��Aq��|�g��?�8�̘
+�z�x�t�ށ/�5}�a��~Y�!O���^�֡��.?��5��#�1��t��!�C?���ې��/�T��T���8�:ֺ?V,��� x�=沑��hG&Do3��N�B.��4L���Σ�V���������v�;��Lx�=�]����	�e	ޙ���/?� ����ChtuA#�$H�ǯ�mʏ�U_J�}�P�;ԅ�����ݠҙ�XhJ�F�9L�����cq�6���gи���y���M��.��<ВЀ�D�5�N׀�{���̲��������S@�	NF��U�v�>ʰs��#X��	f�~���:RF	*�)��DY�������h�sW�T	�p�1'��>Q21��X�V���ib��N9�G��HYW�Є�j�4uͧՂ>
цD�<�$�tAA}��f62	RGPۄ��M�iK���%���B��>���*8��W���
'z�r���Qځ������v��Zb@ٜ��
ˤ4�r��>M] ��=�S��*=t�� Ak��	�u�x�u(M���Q����sx<�~>t�������zl��] ʖ�m�r~����p�l�r�/���:�ʜڿl���k��˾�w�Lđ.S�>��%�(��.}�#����D�s��e��^��I����\�Yz�,��sO#�G�[���[��_PK   �|�X�Ƚ׌  �  /   images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.png�x��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK   {�X��"�IY eY /   images/a366fc27-e5ed-4ac3-9d3c-a6e1ff305d7c.png��e\�-��{p[ ��[ �\	������%��,w����^������ef��7�5]]uΩ�0%i4d"d  �&+#� @�  �lD���������@��!  �J��0<1@� јUw���� �~��A�,炳�W9���O䧂;>���o�~������*�j5#O��y��Zm���|)�i��;��׷�9>�^r����y?������|�
\=����d��ִ�ԇ��Ȍ�l Ix~���6�(``i��@��e�4b�-��\�N��wBS����"D�^���_ku�a�H�c��ΟK�_�wYC�Ѻp���8��& I���5�aǵ{�޴���b��l�/����䍚Ԋ��ޒ�aÖ�¨�w��Ce�R���r�AüE�Wq�������D�L�����mImkI���w����c�}m��à��r��?�;�{~��IRB�'uϔ��4�7��M��+G箷d^&Y;����_&C�'�Vk�4�f��o[q�(E�����5j#��a���ލoI�����jȓJ�	W���k���$F��v�մ���5R魍�˝�\�M�N��VK��+�>��18���Uw�۵�d�f�O�_���<.��k˭G��9�[���w�U�4�ԲM�py��A}�U
?xP��rP�(;p�-J#��銖 �ixLD#=A3~�|C4���j�*!Ǆ#��y���7��v�K�#��G��\���� �4���B�8�A,����R��@�	�<Sj���qW�|���)6��
G�fW�&gL���-/��-M�D4���"�(��@�u�hD#B,�2��F~�-Mo��×}j���n�e��F�
9�y��rPL�"@�*4vO����1�̲)��;9v<��s%�M�|�.�.f�*b��j3���al͋�58�Խh���L.���*�����Q9�S������-�l�t���D��6���.�A,6�����z�_X >j!B��!�Vxܛ�&A��V�ˋ�*V��~U��G��1q��9l�Q�"6.��Xg��_��;�6Ԛ|Jȉ��m�ұ��;�N^?<n�>��&sb���-�����������Iչ?S�=]�V�y�w6�ԍ��(e�d���`��6^%Wo(�]���k�V�E�����E����ңm?��-û#\ٸ �>�}�����q�����/}WxA>ҏQ�~���$9v7��4����D�h{{P�%v�ۿ������o�-k�_�8����<f�h����̶�(}܁ ��$-��#�S/�.w\�way��O�^��Bl���[O=N]��c��?��H�`GͿ�����d�b_m����J3�V�_����1O�%���O��:]>kj����)��	6� 9��h�~�,�~���Խ�q��|m�̙='�T?�-"����dV�-��M�G��,�'�8׊<
-����^�%�	<�V����J��׿�gO������������/r��[U����8�$�cLf{�兒���_$]G@�H:�Gm5\ݜ���
�&*9Ǿݟ��r6�rKu�TNڤ�>�%����jA�\:�������R��Ф�|F��ᝥtx�G0fAo 8�M�����僰_�F��s_�b�Q.�'X-��
������/����E&�,�;��ʀ|����S�ѹٗm��&�I��d�kE{ι%�����*S�|��: �a��O@I�s�s��Sҵv�j��b����O縉�s�\�z���C[�%׊���kL�����������|�%����B��O���d���˰d4�:���⢎R�e�������.�[A"���e��?
��
L��Z�?�{8�����l��%��R<e-�Bu�0���z`~�]b^�E�����vhE��{9�m��y�nϩ%�-���N��y�}C���&�T��ӍBw�*��ȇ�`2�6&H�+Z� y�á����y�"^��e_z����s*k͖��U�5����G'4�NP���L�;�����<֯o������q��W�"Գ�l`O`�G��q�b.����9b�K�zx�]��r��a�V��}Z�z�Զ�ZC_$����f6n�GZa:�9jQ�	�$[�GE}��[�������� f��MRӃ_c?��y`�C� ���/�3�2eg'�Z^���mob�xH��E�WD��3Y��y'�l$1�Z�h�m�4F3G��RQ���OO��u���Y��n/Pl��A�X_H�]�m�����>��?��/@����Z-3P�%�̯uRk�T�H�����P8y`���Ca�[�ZP^~TJ궴�Ǥ}aY��D<o�H���t�nr#1�Q���'�q FRۍ���QX}.>'�g��R��h�)�-^�739��'6_M��
����tjez��`ԡQc 
H)Ň`�k�<�� a��On�D�,������o�^܊8�㈃�#��b��a�k@cї����S������]ZQ�qYڬ�h�u��|�}�~�@[��}iފ,���V�q<�D9L�B�y��D`�#:j�͊�@0���m�ș�.��K�����z1���� z�m��n�b��\�� !_P���aM�)6�!X�pJ�.����{��3n���/ʲE�J�Y��W�_�L�d�h��,O����=��@E��2��h�2{��AקL��V��bf�Z�?��Y�����\�;;J�lw�\�<\ќ�L�+z���0 َ��)��$�S?�n`��lW��m��M���@�g�����f��o;J�6��������5X��뻈���t{�v�p�B��Ll��+7lkD�\O.E?�6��|�a5�dZK������]��@}���EI��/�9qk��N@o�Y$
es��I�+F�����U4K��-	��c�w���~�X�����cM��:��ή
v^>�j"��<�Y:�������l��5,cf-`b��ǭԯk����)ÎM�dZ�F*-{�X@ɹ�Vju�Gg��"˓DU��W�0����k���Y���.������Be�����?:T�O�VI���OOO��������U��.�W�q//
�uu��WTD�t�S�	�����|�eH�s-����/�4��ٽ�V�y����6��c����e�&qt]���xy�%yZN����S��`ՙRC�O�ޟ�ó�C�3���ܾ�Z�Vepۢ�q�"��<RYnUt�ν�v7��u�x.����m�Ε����W;�Ț\���%L�����몫I��z�"�ك�77��(F04p}��Z���}?�ՖX�d��mɉ�*�:�����*�:leאs	�up�5����R��/q��WZ�&��^�\SYUQ!S�h۩SRe=�ۣ�޿���Ȱg��Fۻ�~���l����T��.�5���̧M�v�msZc���7ww�G�Xb�J�r�G��IwK��l �Ӯ�3��('c��F�Q<��(^�ۣ��y��Fk�U�۔�jy�� �X�^��xb���h��"�|������b���9�s����n�fT~yu�U)��5�?(�\}�����RÞo�#m\T����c2�ƟN]ݱC�	��Y7������y������� �
S��RL0
TL!>��6�ɱ�0w�J@l3�in�u>U�4	�A"rwʗ�	�P���ԙ-d��T��/��$|��	��k_>0����_��'�u�'�ؐaZ
Y�ۧ{�3�f��O�M,�k�����8??��Uk����~�gd<z�,E�:�Z������~kV�����%�k�>[��F���¶09JS�@��&W��A����x�2��=z���8�*��8<�Z����7�C��J��%oE0$v!?N�܆���"DtxVw�t��V\�~�z�׿u�����+6|��=Zq��P^\K����>30Q
��F��ۭ��7�I���da-:VG��e-�˒�kv��,��B���}	<�'m�`������)�땏�y^}�:�i�>��?���Z���w�'��#�T7��tT.'�m�O�i������~�Ͽ���ۧ�~ ��2���b �E4��?ؤ���[$�>��#|�d C�w��P K�$��*�s��7�	�._�®��:�0Q�8ax����D�j�*T������!�Ժ��������6�]EE{W���mH��Q 8��F;!�V
�dv�?U��T(�����z���:��3B�d�G5�==I���7j��zK����/�p[��uJj�z��^��d��XdRe�m���J@��a$�7b.�ϑ�!��%/W`Nd��B~]Vշȹp `�����~�`"���)�_O���MF肠�,k�h�a��x`������N�"�+�bΩ
pQ�KR<բ�<��o/��SF���J�X��4-ɍ[�{��A�]?V�0���H����i�4��|����)pY��Q�"703~��\>�/�\NI`d=oa�-OO�F8��t��D�9�<�'S��܆��8y��=�=f�#hy�|M�뮁��k���R�VL7���`lM���}2��!=�n�?��ΜH�繁���2uf�o����$��/eJ�n�!z,v�G0nok� $�ew�c�5#���ikˉ���Ŵ-3I�ihR�h릢Q���%�3`"�B�DD[������a�|T�%r������+W��Wօc@�����8z�N�G��G�**ܡ��.�'��-ϛ�(���d���
�Oo�0�����k��+��8*��e4��nZ	r��a-�T��������{?��z�o�a!��sB`+�|�Z�pů��r�1(*�2n���N�}�W������_�R�q,V���,�R���ItzȠ���]��0Y�*S���hBw�/��|�*sn����y�C����B:�Ym.Ϣ��o�!
MLA鉨�CՆ�L�� X��pۚ �F`�w��06������_�Z:FI�Y謨v�_Y�c��n1��ϡб}b�GĴQ[��~����^���)S����|��/:������q]:� 7*eFD���������<�r
�����v��u[=]hu>X�]i��[���R�q�z�C�����l�����J�<v9��h���@��q��r:���'0mN��ʯq���أL�K��Y)09&G��wd��8�Uw늳0��!bC����)BT+|��u);[�j��1`� ��&tNW�I��62΀��@WEV܈'�d:�b�xּS�$`y�������B�QBj���J�Ť�T�Ч>A}��Ak��>����7,,h£CIg��	���³_��R�06���"�WO�"Ʉ' �$A}��	���\�p��[o	deeƫ�<	W`���##FDM����C���ȏ������wS��s}��Y���z�7��i6g&AYd�	l;�����S)���_��2Ca@��O�Y?���ɸ��ƫ��r��+�)�|��m�~��JG���Ƴ#8�c�{F��h�rܯ��c8�#�k挒�t��$0b\�@�v�����8
.݃�Xwā$��ǋϵ�3�.�L�3�|���]\h���C�(9@�N��n��q��X=d��&�;:��F�V1��u��,��rB�/1�t߾wm����U�(�}��$-坴�jw�pk�Q�J��jl�o��Viяk��$Fxm�M�]�H������r�}Y��oP�G���
��iEjof��'U���[����6¤
ڻ/ (.���W�0X��x����4�	$�IH0��o:Deკ�t��u��%�o+�ԣf��d�(���X+�ˤ��~�<�n�q$?���|��(��^s����Ӳ^�}��o�=��^5v>A�t���F� ���EC� R	���+SZ�"��+�_H�%͢g�@Y�����G�:5�g9�:���k@k��G�:K��.檡��'p���(�pj38辕��J��o�+������������>8�: ���n��=��<�O]�L��}��i0��`~��7���؞�/����چxp�?Zਔ:���� ih+��0I��R@��5K������yɪ]{�3<�f�:KN-s�U������5�r�P���'��ŸhK�i�x�ҹd�>���U�R�g�1�qۦ�i���s����P=�e���c�V�kO�읤FU�w�@�Cڂ�;���!��> ��P��'�"��I�@�<3�JyJ�Q0e!�3��$HD�$L�� ����Y�����(a1���;�Yn�&�A<��^?��]ݦ��,��L=�5�|9ЂOS�#L~АQ%��~-d������C��5F80�`���a끏��핎�W �R�v;��n�^EN�s���Z�����l"L9�9 �,��cWrw]�yk��i���27/��{�H�s�ְ��8_��
1�?+>�Xu����A{s\<��m�|RJShQ2����<ؾ4���
�7A�
���Q���A�YX�P5��Q8���/@Ze___Q&Ǿ��R�C^���RU}�]I�o~ïUC8�p[��"��Rə��N��;8І�郋�,��Sռ{�,��^_D-��$�FU��2�>�����UQ$x�]@�Դ��V��v��bU��#O2�o�����?�j���Q�.$C��l�u��c��7e�|�9�:ϯK���S���AY��
a ȧ�k�Q,c���^�_6��D�����D�f���UPqX`!��1��!jF��yd�T�>�������l1�xy~�~�ە��.�."!��A�ޮ�5�pG�ؒc�7&<��1v���#�4˳�����~_��!��������U@��yT���c��K��,�s� �|�0�{���ֺ���~B?[ȬiS��cҾ��{���� ���75#Ŕ�Ւ�h��HOq8ڴ�Y���5�5?A��xS+�5�1��<���9�O�gW����r]'E#x���c͡a֨����Y��E$�;L��e����eꙛ|��L�p�/���F�Ij��ڝY����d���(>ٖ�����(���3�?C��?cr�2p��H�m.v_���7�y.[w�����˺���gw4�u��������W�a�Tq~�`���y�%�0��	l��5d�����Ǆv�/�f+,�>vf�i�BW�!�Φ��V����@pK����a����P���(�h�c��,��A�L�)�mε��<nKU��>��訍�(�3�=Dp��Z�F����z>K��0�Ц��L ��Q���-WCug�B�y ��rt��j�bmqh�#��U�h�*�oo7�������mΣ�G��qJ�u:�N��v�L2��	6{���il���:�t�?�c&LS�
#(���9�׮:R+�j� "푯��&s��2�O{#�}g
e�|�36^�ls��ը6&Xk��"[��Ğ�]@��C_(��M!#l���L:N:��I�զv+��9sSMwޮJ>�k@�"4nE����]���4�f�Z�&og~����;��!J�W�خ�|��[��@ ����+F�����nJ��`�<�a�rm�3 ��J�ޮ��>J
��)$y�a�ǩ�s����ؤѭ_�Y׼ţ��b����S�VMlU��ʲֳ#Y��|�$�d�n��bj>�VS��K� #�?����%N��+�����)V+$�R�5������]�������,�W{������G�"��u~�����5��*񐲡���=b��j;N�:�#$	��֋�G��!!�9�Z�Y n�`ic$�r�܉��p�D���(������G|�6�KJI��edI�^A�4�|�i2������jI6��;���c4z�3>Q��+s�/��Q>�a]����T��FT��+$���F����&m�1�U���ٯ^g����Tc0s.�۹[���X���}[̹�@=�/�^L�.�sW� q� ���6�2�P b�|�������`����{�j��2L����T1���c��ߞ"��n��}��,��Q�b����UC�A���z�H� ֊����me#��	����P�Χ��E���
��A��t6e\L��h��:h�Ԅ�P���N 	�$��#z(�m,X��ͤ��J����x>�
%���K1z�H����~`1����=�Kȼ?����?-r"��x���En���8'EG�Z�������{�K,�6����aƨ���3ڥ���6~�����T��rT1
s���l��6)��I�q,���*Ċ�WZ�$����~�T@�ڷTs���~�X�k+���`S4�kϚo #I;r�iV�~ޕa�����
FàG�c_\j��F�!�_�Wt�U�1��c�?����KZ��ᴦ�u�p�9�r�f}/��d�3�$����J%����e�+��?tE��V膇����x�a �@*ꈌ�R^C��ݖ���h�։u�����;��c
]5ARD@!��<����u��<Py�m�u�ά@,a�X9�7�������w�E�?��xf�\��1?��vX�P�V=�K�܍�kN���Ӄ0���L��.�1j"���lvJc˖�"�%X�>�~;3�f>��.�+��Q��5���u�h�ӷ���PL��g\F�L�e�Q#'}�界ru��X�jn�Tac=hw�o��g�Ii�
ì�L���ўK0�$@o�������X�#�K
����e���C�B�=�H�M�ύ~A���ym�b0o��*�i�(�K�1ӊ��������U�/~ͼ8�/�?ԓv��Rם�u���w!O��*ΝM��p��⭮�靔���?�Iq��N��\Mŧ������6�O��q�a������`�|��:��tVi@�+�HI �s�)�˘F�{2
$�lE��Q1�\\}�e[ۢsv�N�ug,��(�T��
�i�ޯ��Z8"���G�9�������m� ���-�g����llV>��U��E��x4����Aq37��D~P�پc��^��v�֦�\��u�`"�>�Ľ67�o	�j>��t�[0⃡�d����8'_F2���*o��B'��npX���eٝ���|b���l�7O����ҰY��3���e\����aԗ��<' �}�$>�9�Ͱ�����Ԍ��FDD.I���jo���B`�ˁ!|������^F/#`O��.f�LCwr��t�#�Ӄ���O���Yq�vK�crI��}���l�:���NEv6�,M�ǻ���*��fb}�0L����V�	^���yu�&���g�!����������$	��Ws��|�Q��|���p��[E�@X����?6�c��3����Z�������nO�/4w�$.�d��ג�p�9�⩛5�"�4apo�ఔ`�	4�cJm���?==�(��%R��ҾO���k� w$n{^�H��c�R}�Ȅy�9�5��j�UBs'/Čb�\-}��|���ً�*Ϛڱ�y
8�06��,;�EW���d�[�~�����.����b��^��b��{�;�X9���d;ޝ�V#�(���UxF�C�N�ǂH��ʵ�o����\���2+��ջj����|�닞¬Ь#�D6<��i����b�ϋ��e~fWsQ��K��\3KK�j��m�04�H�	���].U�v�m_��JK����b9#dPi��9CԴ�^_E��Q�ժ^���tdG�w�hp]��bs�lѦBU��)��>�C:��U�;Ξ�YWw���گC�phёO�ˋ�~�(+O"���誫�|�!�+�p��y�GyT��/����^u�l���l8��Q�˓������{�C��\$�M����`,3l���	��Ήv�엻m��P��KE��*�h�*���`�����(j��)(�kK��kMc�-�<�_�c����F�e�-�;�E��N��Hٷ�#K./����7�����!g� T豟��]�4���m.���%������֐}/���=��*Y~q�<�Xu���gE�Bu���(C���Y+!o��������sSz���+��a��ٲx;,�@3G�r��^{\u7��n�4��""X����V�pd3Ič�!r0p�+S�綘�<'w�7/RP�St#9(^XX�8�7��b��k��naZ���^�ZKa�
�hhEA����'����J��`pB;�B�\FY@�����翄c��s�۔ظ�p1����Y�&�o]\��h�6K_�S&ĸ����Þ�� �xqE��z���l>mҵ��q����P�������+++�J��7��ө�j�}-,n4~k��N�m�d[cC���3>U����Ku�]����L ���h�\���jݾ��i�E�+�6�7�dH�=���#tJϽ4�yL,X�N��|�K0a�1)F��ql���M#Q�YhsԨbkC�F����t�W�l~�UM뺡�f������F���ea�m�Ŕ(�F�g�]�7F[q`(5%b�]0Ůu�C���At}��Ԅ�BмM `$���O,��R�n��)<��F�^��1BWC���'���v�Ĳ/�W[��~k�ʬ9�Ԯp��3e)-%�Uh">�]�!���|e�J/w�`��%��*��p���g>�j;�!%M)̄uh#3ޡT��1VF}�ko�@��-���w��w�$�d�|�xS۾Z�QJ�B2�0P_�`�U����g�Np�����7b��7��y]#���/�4wޭ%�(�_O6�rs�Fr�o�ttN|�%�f�קb-#_��r�����%.��r��Mg�~�G8��)�ܒR��V1��{cҤ$�\G��ߛt��رg����f��%R��*J�[�fY�i�`�A3ԤN�f�
k���N7�ߣ�@�]&�-�^ɮ����^�ֲO(/��	���"�%��y�:�6����C�v+��k�wȴ�3��iM�������b��S�*���*<�j��b��V[\\��-������#[k�o�$%�@�����;�Y���ş��N�Yd��/��l��@�@��ގ0N�>3̻@m�ņ!����]�֐9C����B�P�7��C)�+��&��p�l=�\��:B��p��/�|���[_l]{6��L�B�C����W���?0�eWz�\t��8�/]�eC�t$Y�cz�����D���7sUo��|��:�2��@2��������wל@�1'ܯ$lK�����4�$`ocߌ�!6�di����"�E,C��s����^�@�;�m=�~b9��3�w�i�)m�#3�Nu@�����u@N��V�KcO{��+�<��#|�p��ܱm�%�~�Q��.9ܑE{=ɽvq��4��ց�#�P�X����vaF�u8�����J;�Mk{YDȕ�{��P�JC���L SX0�P��`�����G\4.���A��U)7(�9c~Vy5�h�4�+�'��M9ZWz��Ԍ���A_�����*�6�a�$Jj�� ߘv��.�����`]�Ѐ<k�J�������V@v8��X�c9���`M'���A=��ں`BKH�e/`�d�]0k�����S�hZr���`�����R%ȁg���B��Tl�$n�������K�@�rߍ�n�Y�����ɶ0�LA�I~pe^�Bw�I�ZG'�'�0H0��:�N5�u�Jh	�Ĩ��5�c3���M��lL��=�[�MY`�����q���gDu��p�A1��:S��2�|"z�4ݦ���ɘ/��,�Ҩ4�%t���S�$�LO�Q>B3�NL��2_;U����=7֞������&/���i9U�a�x������"8�Foc�caEޠ�i�
X�a�v�x�]����O�5g~1�i�+�zk����FD��r�qD����p3���i^��N����� �����&�S��[n�S5�H�5ĒJ;+�"� ��g�����B��荋x�?��J�bC׋P�+�o�#c]!n"\
Kɚ�T�
�6�i�3��p�\}�פ�a���O��Ltg�D���-ͨ��w�,���2�W���P~j��$�N�vsu�PpN▹�PO-l(G�Ƿ��r��mQf�a�=]C��_$4&1�� �Dܨ�(qqѸ~�)��:0���E$��ZK�����|LL�}&@ս<?����+���?��A�|
Ke�):�O�c7_ ƹ�x;��4�� �BĞ�t��?���]M]�����/ bs��O8�����5�P���J��GnifY!���j!&"zr�&�5�<=�Ԃ�
�ISx������pa&�G������
uGG��	Zv�����ȳ�*�^��RB�Z�.�j�D��f�n	F!1�֝�3e���@VK�Dێ�Bl �@��^h�ց	��fw�bJ�4.��晌p����ٷr4jm�{��('�'�7���@��G°��Z��q+ip����%����Lm^� 1��ZDQO$"/���(΂��j�.d%@�aW���8��Y��v.��Kc�����>.�g�ܐ=�ְ�����&��5\k�
��}^�szB�9�P�UK��t4�s�����c8xg���RX̰�3X~���o�\[��ԶT�v����y�t�y��;�5�1b(G(�mB��K�7x�c/�X����ʎUP�++%l�|�NҨH8َ/Aǫ��~��e��H�,�A�׽�i�#J1�C$2�,$+�Q�@������T':V����$R�tZ����yђ,���Ԟԟ���|�c������'���F�{�wk���7�#�5 ���Gb3����i�DbwG��v_��~FI��TlߜA#�`ґ	��A�IҎ�3���O(��]'!p���g� "U�`1\�P��eu�	m�F�~�ʨ�;Z��vDG��B�޳"�ˀ ����E��4�_��U1�o~��65���{u�E��]�8�HD~��<�����oGycm�2�?9�!B�k����%6�,,h���8�?L�ZB9��ؽ�z�I����|0�j~��ށ:�TjR2ѽwR ��(��bր6�X��TD^;�Q S�V�i�V���~��l	�C�@�>~��Ȁ�қ�uDo:M��V��+�SKL��a��l�hQ9狅<��x�)8��d3�XXrhY�G���%��[֢�G�F���"�t�ON��)�S�5sX��db컗�������|��ɔ�����59�ސ�b�HJ�4�*Ej<���r��:���:��Vr�)F~i��q\u�F+��s�_�/�rN��U���K2'��2��������.�N�"���;��U�
%��T��v,�}�i&)n[�o7%��2A����r���#�P#���}h��4�%���'��P)��)p��@�Ts#�^8�st^��Z�����)�CE_u�J��E?�+cDTJc�QO4
�-����w��,T�2�;��R<���;W��/o����"�e��Ʉ?=t� '�SH:�O1��pjK��L��P�ۣ	eCI2�2��w�$�6â�T�H�cB��O�j���X�>���S����f0���sh���7���	��;���(5���?���/���3�ny��_σ,��4��
���׻eN)��3�6����n��ARw�����H�I�w� V?�4qJGI���SZ�T���������m�O�J����W{���<�+�<�C�?t�Z�AIA�3� 6�����PRb��C��j�W3� կ"a[}�lLKl75�'?��Y��u7w���;�}m��fy_��i�P��3AwH��/��Fw����18��C/zyX�u� � ��c�@���¼�E��ge_)�5���>�@ �a�%?��<��!�8	ikcc�Ņ�_Z�V*���:c��@�އ�4�A�D��%-!U`G	Zw���Y�I����8Y���3���p���!�,�T��獛�>�z�R��0��D���FN�����l>GJ�_��?�n
�kY
�5��|O-)~���!�7}C��HD��0��q1>��I�+�!�Yl����,���LMƭ��8�Bq�Lxb�L����]ꐕφ���|q��'��S{�c�P�׿�����EEu���8v�z�Ν�9�����Lς�_����ȝ7W(nC�z�����.�� �8l`
����yw�4�2k�P�NQQq,��
�����#-G����� �[�3���\�Ԋ�/2����c��gp�>�V����]@�
A�#A	�����^g�Y�-���F�Ʒ���GrlyC�!6���U_��`���Mafm:3��*o�܁����v��q8�����yVV35�}}��Wڢ]���S�����P�x0
r����~�ҍٔ���+� `K=�x�[p���Bz]�x�@�d�V �! �M�	��X���n͈i���A���E6�-�a"pH���cGB���1���L (�@
DS�.��t�Bt��5u������h�ll@z��;�h�����d�Z�_Ƅ��0�t��?ȁIWQ0�l�a�J���.�*�%���Hl0q���
�����!�Uua��S\��сDJ�����	?�&
a��t��n�No�y�<"$) �&��~	�.�ͧ:�	�f,�]�旇�Ů;�豶���z˸O�*���EG���?m����Pb���ƣz��<�� w=�BҒڀj��c#u{H�
��K��(Ky�)�6{(ߖl6dO1K(���d6f�|�>��r�e� ���B�}��4&��ڃ�4X[o1�w��g�.�A-�0Lh���<�*��4,"�y���'Ii1���-��蚶1�����F���]���I�W�]|E�0�{�dM��ᶡ6�������������~�$d0�����D8W"%b��[�R���3��|�ؽ�IM�6� Ɂ����aۼH�Ze�ؾ#.N�����f�@���r��s�
�hd(����Io�j<���zH֛�z@�ɩ����_�uE*�'�V�ap����h��;�~c�(���!�M)Oi�)gt�]Lxg��	���#��g�0��B��v@*f���0�,  �K���J{9J��p;��ì	�_�y#�@*���~�i]s4���Eh�����z���{��'��ݗ�����J �s�+�����$\sR���*���p������Y�0���d�,>��i����~�ڼ�'��=��0R��1�,��I`'�#f�`��CUj�S^���D�;M$4}���y�<��0�48����L���M�qb�����BJAQ[���a�4T�h@���e����Y嗄�J{��+�i9�%�ǢϺ_R>c�A�$ @�P0A�#�����s���vr6l�HPFP�i�2̸`�@�I:F�-J]-8�^�h�?a1�n�)�fX)
��5�y��UD�t��@< t��e�悙�/��n��i���@����������i��ԡl �?��BZ�mB���v�~xMDے�3|Є��;S���`���	�z>Ø��KK�ٲr�'Y�k�[`!t�ųK�P<��zK��:m㞛�0@���EMN?$����}�A(�V�����F��C�I"���BC{��$R��KQ�$�?��?�N|����xC=���ql���F�]f�tK������ֿE�9ת�Ϝ��T�i[Ռ�����|��٨gU��+��@ZV���Ģ֧�LN�fY��'�sSvmZ�q���Zҍ��!mx�w�!0���3�DGr�(d��(q[��,�ַ�Cd �2%�p�A���\5H���ZY1�l���Xڌ*t�*��;<��SH�j<�+o}���Mk�ە�1�N���xe�G%t�kk"�ՀSr��y�B�kίt�_$��oZ�T���2eG3X)~������84FL�k��o�-��wI5�d2��jB�g� j)����/"�kS�8	�UА�kbZ�K6D�ǏZu�H�\�hc�ɶ�8�p�}��G|)d�t*Ȝ�=q�'�yy�0��t��
�p��*�)A,�E!)�[�w@Bay^����$��we8V����B�\-� r��,!��>cH8M��o�)�*�4���8UJ���"����>���������`*��p��{�n�h]Fg��0T�3d�f[r�*"��.�r_���iF<�̼3����ƆN�p�������N9ݸ��ք�nI�2h����&~7�~�e)Q'�����{�Z�a.J}WʉB9���N�-��v��of��.�\���U6L�=�Y@�7�	杀�s�Uw6-ƽ%�4���@t���� �t���v`����A����h;X� '�,�B�E_���+iC�� Q֖-[�q"���f�w�}7�ꭈ���]zŒ�+
�3�Z0��c�m���)�!�2)jUs�>zu�˴j�f������B��*�'�d��� ���B�n"ɚE�=��ә�/]��c�/��b^#m��<4@Xw����X�,���*E���v¥tՁρ��'��`��e���[�lP�����h�޸� ��6@���qV�KX	j�����p"I����]��oo�9K�n���҇�p�g�r��C sbvG������h� k l�"�J��o����"���z�N1(��g?�g��فo�n钥�Ϙ1���-�Od�@��}�m�N��a�9�DGqgQ{��g8�/q�ೞ�Lt�=��eˠ����y9�H���̝;�Se"���{.� @C���+3���Id�Jh¢/sSv}����8��4��+���� �C�âYn�?��]���X"�$*"�� ��c��At�_;���* �&v*GG��L�P�&Gl�Xad���^����_� ��!C����f���������d`��X�^�#�Iރr {B���7�#m	�Z~�u���(�Ţ�@ =fi"���K����ԔT:� l��_�}���~�#,G@@���`1��*2��5��P _��H U�.p��1DO��'>A31�3v���B\_"���9܏�2��rHY��p9@��\記YAzB[@�]��tNY]��㡝���@��"3$ee�r�p%�D#�L�P�=��,G �����Ѹo���� ��� Z�'�p���>e���.��#���o��wQ?�I��aQ�,�A�(��K������Da�N!k.���������*΄k����Q%�����'��\O�>���4��;DlLD�C�d�PD�����
d���0�E�
Tc* �y#F=LM�^R��K�!t����ߩU^8�_���ԡ����ld;8��\>���%�\�!CX*�����}��%K���mRd�9��) 3�E|�S����v�1��M�N;���c��Vr�UU�q��X,�5���;bW�Ry�GÇ��XĦ��ZY�p��/D�\�n���|�v�,�3X���e¨�,�3�=H�'�fx�,���5D6�mao��F��xa�1�	x�&˜���%U%�@�8� g J����T ��~ɒ%�DnP�)h8�ԝC����TO�>��< � b +��#@�
"
�a!0���`�0��V}z �Tp>K�K�'��e|�녕��(���'��@���_�2;D���_���R�B�B�<����z4ˠn`�f��lS)��^ �x����\���� ə��y��S��0��<��nm#��`�g��r�,[�凫Yjǖ#`GHP.�.fݲ�	��N����-ā+�D��, ?p�a93��s�B$S�/�؆t� o\C4gd��k�Zok��40av�%�y�V�!�l�Lp���P�9��	���'�S�0D��Y��\���7�'(+�D��C&\N߶���YйY�i�$�Ơ��^��e�{Ǉ��$�Ph��b t��:t]]��t�eG�[��ާ�XE_q]$ٲ�g����6�+���>�H����O���d2"ݫ\&,˖/��"����&��>ș���(	Y����I��y�x%۱	pd�W��C�Ůz����f��ZZZ�U\�hغd�H��I����Y�P�*B[;��0�3AR�Ĩ� !��tS�o�ы!�x���YY'M Y�3*SOa��T����5ϰ�\�g%�@Xr�~�_�A���$��`��uG�����>g���*�L0d?�]7�0���`��o��rx��͡T:N;��T"�æt�#�Y���#��K��]�i�0�> [w��e|q�-9" ��p,�?(��^@%O��6���r��cP�h��%p
3v����I�Eڧ�ƀ	?���rn�AxX��R��јͫ|ȵ����8!vLX"$� F,�	�a��sNd97�w[�P¸zܱhi�����0�$�A���=���mu��5�\���!RF�@tJL+1E��/t8	���<W��\=��l2<8�l������C��R"�A5�1���7�ܴq+�{]��j +�D��^��v�A�|-&%S��{i�^�s?{�u�ԒR"%G��GV��Yl*� ��ñ��U.��LGw��;y���`�K"/q��;!�%�j� �=|���`-��6ᆭ�~��`�X1��fN��]�og\=c:� �taǨ n�Gc]L��ٌX:*�?��;CdU6C�u�P���U�r�0�10"#���zv�bօxqL)!Q@'�|"��s�� �@���A�lbׅ$Y�C��9���h��u��h�ȱԶ����p��jK�l+F�T�b1�J��uS]}Ŧ��9��Z�#5�x�J02���1���3�z/��+�T�!2c��U�F��p��X�N��	~H�S�9�1r� �����B$�,۶��dɒs*΄�un�d,�H&�,G�1T��e���,�+��l]W��eDp��	�ʻ[��u�2V,���2��v�J�V��<���s���:��О�1 #h^��Ndv%��ۯ,��)�) a���L0�%R�t����9��葿���珔L�����*��cQuM�z{6Pu�G��z���C(ѓ�_��z��)�Ĕ��L��uc2Dď�U�����aܕ�`�~�w�ل��	�$4ъe���
ڣ8NESFy:�	��H0a˲lii9�� �sЄe�\Ĭ�c�;N���=�~C��
��8.���d�:�fK0����G/`L�WʔN���!j�,��rv�֡i���Rs��<{�ˬ �UO���"4�B����5�j�אَA��ɁT���>���2S»�1�.��:���9��mS7]��[����J�]1�u��^&��&Ǎ�at�QG͢�.?���g<|���t٥Ki����%��5̂�b� <��S]����aѢ@�\E��6+��ܩ/�2(69^pI�7i���l�I�H��1:f	��94 �V�q�����2�z��{���%2�	x
��ߗ��) ,[���6)�(z��ש������ib�U�4ȕ�`�|���.��v:7Tv�Q���\�$SNc����k�ԇW����g¶��pH=Df͘�}�������"v����?�-]s�w�Pu�Jۈ��{��ldQr���I�g>�x�}�Ewu�袋��G}���*r=�c��k,J$�X��\YP��d�:���-s?F�%�q�m�䵰L�0a/�����#����I����t�@'f:��g�l9R��e�축M���qKȂeY�x�p!���B�uM&�u �6�_#��} ��ʕ�Qo'Bf����=�Q,�_i�r&#)����B��v�w�E����g����R���5�G�̚ <�H���{�5��X�%:`�T�x�G_��{tǏ~C�UM����2c̮���6-���L�5)�s�1�ŋ΢Q��y]��6:����Օ�ɠ:R^�#"��lJ�:��[p(��_1������:�LT�U�~�1��YO��@X>}�\,�N��H��8儹��>;�{ ���/^|vESY"w��0{��ݖ� ��;�@��]�{[0�� ��gJ������Jf�1И�V��#��Y@c���Y�0!�	�����~���e����2�DF��ش�t�Q�i���я?���wQ�WQڱ�@�Z9@��z=�϶�]<����(}���c��x<A���~�ӟ�A�=Y��p�CZt�-�y����g* (���
fFy (H�3�~ f����'�}�, ,�$�o1=#Ć��f�2��R��yB:���+V�8g���{��{ʐ�|#�e��[%�/�T�NF��Jv��F*��a
MES�Ҏ��Q �W����Lt$A��N^�������X�Ɯ��}�Di7����lJ���o��1C�l#�d$)Z�rV��fq��$UW5Q�!rU�s:}��̣����j��t���"��ck�{��0�V�����+G9�g�Ad������* ,�vp��������a�f��'�E$	;��q:���H�l��� �ͪ�m2��
�n����Tt�� ��	O&�°��̒�d�w	�ֽ���v�L�C�꥕+_���8Y`% 1�,8�����<��������_C���҅��4t�8:�������(ք���jiJ�{��;� �I���y����$�4�B�
��;m��! ���]�E� ��C��R2��H,ʻ��%ۈP:��6�Mv����7KLK|b��>�zM�x������;Fk�;�d���S�r������W^ynEA��7j_wkM�{��ә���+�k��#t�~� ���5�	��p�Au���/Ȏ�i<� c�x*�dv�:�7TQ�LJ_-���1�c�Ow��|�^x��`��SQ<��a�r�}@�1�2Ps�4��v��C��I���"� ��ҞK�!�b�h���`��b�����qd9�0�8���L����e�BLX|Stv[�g�.e�\	]�5
�lXo,�dS'�Ax��˖-;w��魃id7�l��zk��5)WtxBu�蚯1��M��5���ܱ�L�|�U��a�r�,���o��+�tI�h�.�a������������
u��N������c1*Ή{�巍~P�m�
��Kv/��f6��������X�gY1�OCԂ5)����Nd������M������0_t �2扦��]a����ئ�{���yf:�f��0a=�ד��L�	���g�BW�w |߲e��ms��Bn�	���N��BŰrl@��)4-�A�s�lp�Ż���� ����~4d���ӊ`�r^�����TXm�r��^87{:�w����6�p�	 �~���ֶ���@��ة�8]�gb`��5�6��$"˦X,B���c>��
̖#5�\_�,$G�kC a>L��$yn��qҰ���Vˢ���F�r�9+d��%s<��[����z��dG� ��,Y�+�rQ`�����I�2��\�U�aܷ|���*�[Zo�IuMB��D<E�U���dG���rF2L9��	�e��$UF�4�lBJ8$F�)�>�隱x�рa(�=�~���2U	kʌȈ���#�wf?�	���ʡd*NQ+ʫ9~ҴȴmjVG�M1\^��0_������`��{$���З,�o[#nu�Y�A��+�-^�'Y��%xj8�1(+���[�`Ov�0�o}�^la�Ul��>#	�		��|�6�%׍S�mQ$bR:��^�8���f�u��B�j^y��yWt7�I���ό��"�r= K��VObf�|��ÑL��,�@�� �x��">�qQV^�~������G��xG��>;g���)��m��.^����3g�L��/G|���M[Zo�%:&!cF��H-�`}M��{:9���C*K ��X�1x8�I<DT@e��ȳ�>�ɑ%яhf"����908�(�
�8O O@X���Y�Z7����]���R*N6�$�IɄK��"v��$�	"�!;
	1j&)ׯ���GG��<����;63ʹɧ���{aq�	 �^�&,;x� ��b�Z�[3�
�w7�zup�{�I�`��L�ӎ�d�d" $n��V��Ӧ��CS�΢�j��E�[�|v�T�([v�f���|���g�������I��?��o�C������f���M�G��yG ��4Y���Y:� l��T��)9,p���x�eݳd	�\Yn���͵i?w����1��������Q�|C:9��|"x�Rا	,�Ǳ�',T�	�׳a	`JN
+��4}��.��z0v6 ��� ����Z[_&�H��ɱH�5���SQr�AV���a6��4��5���;��wH�[by�Aٻ��e��LA��_�`c�`߷PފK	��[a�,�>�Uib� ���-XĤ
$�6* ̣M��/X��*�T
kO)j�4���jklNs���U�`󇣨y�Nd�H(�o��,Iؑeq��
 ��aGu� F=l3����^z)��u�]�dO�S�Dx������ ��^�L��^a
d�Cy�+�c/L�+;6k$ϳm��ŋ_0k֬u�i�E8�޺��LO�TrrG $�����9���7��-F	<��p]�Qd��4 I�![@w������h?�F\5�s` �k��H�P�����w�R0:���^��Y�G)J���ݽ�b1?�r�dU��[hŊ��֭.ّ*�.Ǔqf�G~�=a
��.��ϻ�`���X�B��̪ �U��g�@F(��} �K�g�jx	(@X��更����a�ʻXD�ʤ�S`�!>���Ѻ��ɶS4���>�S�}G�1� �xJQ]�pRf-��DK�UWײ��Na[���i�O~�LĂ�q�㫯��������9s氜�裏���!���?�C��ȓ�2������%��ʲ;������������>C���D~�hѢ���-grOo3a�0nn��It���M��x�Lx2���3B �� %F�5��7��'d��p�@�R��5���������>%Oh ��K"��@��������˒D�;�V��$iܞ�����s3E#u����􉏟O7C��%G�)4g�?�|�(���������Je�ʻ�T�	�re#�j�GH�~N8D++�`�>ɏK���m�4��0�a` @�[��6/ۊ���Nx������G"�륆Z�/�O��9��V�����^j�HS<aP4�@N��>S��z1��� ���G�!|o���1c��y���/2�A������П����7�̒����@`
��P�ꃄ�M�I$P�_�XX|Z�C� ���{�e�����"���-Z��� N��z/>L8��s �O��#�|�?|c�#��9�0ȊC p�]5*��[��Q놁q�:�(:묳x1��s��N6�mI�%+\p.v�����7�N�����:=����F�l�̙{�n���xo�^}i}�c��4���(�d�s��t���e�roO�L�����!�����E.����Y�pL�9����|W�����;����;��Z3��E�E���g>��O���sB�P�+_�_���DnE�]�x>�|ұd��J�ko��g�}�&�=�jFS*aR4VO�
R��sv�0������a	�����?�����3����d�©��������'^ G`ta`
�駟�~l
&,a�����*�u���E��p�������.���-J) �p�*
��˖�	E<"v-��1��<���]�7��Q�b�|������x���l�=�k.�M��\0�O<��xE/��B�
]u�Ulp_���������׼�y�vut��W�ڶ�@sN=�.��T��W^�Dg�u)�kMYu���r��� M����^-�(�����s�����Lh���\c _�/k �K��cy�r�+.3���}5�c8���� {����L��,l 8�;���;n%�레�K�z!���㑏����7�u��]���i��#(��)��D5{^�}*�YL��3 m���C��R�8�́�b��~.�
�|��\�8F�_    IDAT,��<��.B�d����?:�.A�����cG�O�m۾kѢE_�(O9w����kni��T��g1���/Pm]�|������Bb�͊sM �����(�P�d���=v^�f}�H�y晬A��/}�G(� c��C�\�&�r$װ��E�o:�����詧�JӦ��o|s�3~z�����ͣT���	?�
�W`���79����Qc������k�>��+K9V��a@v�eÅk��8�xa}1�3�%E��tr�i9@8��JU�-^|}��'RWw;-�j=���4z��w��4}�!�(Faf重b"�%�����u���>��>�Cd�������±���+H��ԧ�3H�
 �z����(�ɕ�<�(.�!�\lf��������g�毮����}ϙ?s��ͷEz�L�i~�F���g�m�z��'�̎�_q�nZ�P���#`D��3k�,�X 3�%�~�1��7�J��r
_���cP���Q�!1J�%�a3?8���*<iX�����+_Fo��53i�U���L�Wm���9�M 8J
��(F���~���AKB�B .��#����9����b��$1��Co)=����	0�Y��~��[(�襆FE�_�Y:�#�Gt��W�SO�Ұa{З._D�L��'�1���Xq���L;���J���z��N:�N:�L��K/�Dw�qmذ�/^̑7�x#/�8�/q��%��AV=��2�H_��@��������~0H��tJVṑ����._1��ɓ�Ʀy�#&ͻx������${�q�]e��	��=�^~�Ez��g	���� ¸A	'��1�'`(h7�
��2�
`��a��g�i����aA�q<>ñ-Z��� �qMLAp���>�������t啋�����A�^��&Mއ�{�u��GϦD2Fi7J�YEdD��9gp��q!���Ǿ�,  �曯����	�vwSuU�/9�N��<K����7��'��iͿ�2�c�=��7ͬ��N��㽝��C�����А�v/^������s��	'��}��?�}���e���׿��H��={�l:��=��;^� 	Y���υ܀������G�����M]��
Ѝؑ_/Z���Lx�s/�6r�[�ե�3"xISt�!G�	'|�{��f�2]dK�%��������L��w=='�PBBB "Hii�@��҂!�8���w����f�$� ���)�؝QQ�+�9m������OǓĐ'�u�u��������_�~����?DfI'Wp.L�����Z���p�҆��68���"|���P��r̄�6\�n����^��]{�n���q�����[�ՕU��R/��1��� L����,C}��%�9�t�}�*�rjk-k��߫/:5�y��g5��V�Ԫ[n�Co=��`�V��4�<M%��7��d�~����[�DE��6��;묳�S�����'�ֹ�q��8�Xm�|7������8�b�s-�n��N}���3�ל�r7o
�S�V+�T��;�ν���L�8���=fӚ�z:�F.: |��O�y�[?��g�a��s��7AB��:�!�r!�)��@]��Þ�|�K_
�{��;<��0e p^N'�fr8�c�%�s1~�bHV��ٮ�������Z��I����ڔϕ�nMY�w�r���%Ӥ �f�$O~G�?�����k[�e+���^j�&}����E���Ƥr��^zq�~�����7M��_?��_���l0fHS���A�!l��	����)G�ڈ#�y�����?�A0G��7q�y���d			"�t YH#�P���+w�h�r79`���4L��JWM�SO�}�]7�r�)�WE��o9j�����Ӽu�1�1�2�������^�Z*�IPI� ��TX;�� k5�5�����Yp�q@�^y��9���<,+戾��t�؎5��Љ1�=!$-�}�7YU�	�Sz�!l	�U���P�{�K��1�C��ɪTM)�	��4y�t5n���!~m��P��FᕫW�Ա�CMMe�}��5mƹJ���Jjn��[Kڴ9�|>�Lj��R�{�q���tD/%���1�Ad�=��}�X�17`�%�!�c��v�i�q���6��"�O�+����X�ҥ�}>8���Y�|ꩧ�y�ۄ��L���wr��Q��lZ����?��,"	^�a���ks�F}���U[#��W�X\p�/�a�e�sh �EP� :��dђt�+B�q�� 1��s���}��� �j�☳(�����\k���y��[3*��)��kX�H�������ھ����&>��*T�԰W	����vH�	0��s���@�ZHh̨V]u��z׻NR6[V:ԆH�\kTwgM�T����*�Jg*a�Ѱyp*�+~��<�i��aj�[�xm9A�7���G bS�N 68;�u�ĉ/���f�,0	��h�+�=�F�tWOwg2٧�y���0~Ӗ�����yՂ���I�#�Lވ��:u�8t����3*vcG��h,����߀'�^<������9��H?�&��q�{�F�5? 3�����/� ��a���X�`SvP��s�)�8kz��O�k���BO��P�2���k�(E�rج$N��K.�l��UO���x���P;C�/��C=��m�n7ftV�U��[�m�*U���ǝ�7��r� ���BoAz�I�,[�kD0�K���#����B�0���ի��;��N���I<'	Q����w`��8��`����ӟ�e���V�@��s�D�Z%c�s�����xío�i���|׉�d-I-��d���Stҩ'襥��r�������z��:i2:	���Fh/����C��6`�>���SO���]�Vs��	6c��m|7(�F��6M&�N���gU��:gRd�P!��>U�V�V�as�ƍW6C�r�@�Ƽ��kH�%+i���Tʥ�%ns�fʪVzTKBrjjl����Xe�#U-g��ܤ���`��ը�V�K�
[454(�ӼP 8�$���2�!V�����,=a�u�5��H����P�j,�v���k+v�&Rۃ�@���.����j�J)˯͙3gp����_^�pT�<�;ߝhmjU�3�7����2���5��g�5k��ES�ދ 錗f� "��I�-i��	=���3_(ڇf��@TT"`��k,���7�d ��q�۵t�":+��m-( )_`Ś��F���QBS���QGMP:�[����~!�PS�Z1�KOH�FU�Ez�N������6��Qo����ViPKK�����j���z�p>` ;��9	V�z��a��s��F[�3�ӎ�]̙�� v��6mڴ�z&��2�{�F6��ɢ�j���}Y�qސ�k�H���ܹs?4�E��ћ6,l��6)�I&��/Sa��u�X������MZ�|e�`�m:�"�N�0��d�j��x�t1�`r�Y�pZ{?h6�f�-溸� �����v����^\[��|O=�;Ö0�P*�6B�Wo��a[���
A���Pt�^����$`^�v�>���T쪅H���4jX�O�Jgq�Q$�Qg��B�:�ڢR� %;��)U*�@��G# ��w0�����vK�-���~�^"�LxhBÆ�]w��#��v];��@���8���xa���MM ��G[Q�"HP @�v���Lx�A���ͫ4to?���A����2h��*��:�Lw�[C��@��8:�Tm^���/t��? ��cE=���P%��% ��DG`~`9�&ta��"��7�!8�=x��xƌ5�(�R&�m���eU,oWKKB�JR�}~�>��g�eK�������Sg��!~���P�Q�+����ROU�nӬ+/�9�P�,�*�H�FU����u�R���������p?Ha_(>0Z�����?���%�)�6u�z�Hڊx^�s/g�b����Ŧ��z�OT��8�_	_m��QZ�M�6q�������	£6�Z�Z�91�N$�@��F1���+ۘљg���?!�V� 1�s99k�g9�ҀNq&�t �������\G�������;��@��a�$k��w0�2ib
z�ڵe�
e(�פ�/n��ݤ��ʵ�  L���(C�A��C���%�	c��֥�6��;ޫ����/D���`utI��P�I�r���l�`Xg�;|*.��5~3���RO|3���0��~z��:m��!8�� ��?f��W↹ ��~��6 �	��b� ��x�z�Q@�����Y�R�>��J�mI�=eU�5�(W�Ѱ�vM�0Qd�'L� G~��� a�t����g{@�(qu&�
"h�9;��N:�t���(�	;N8~}�a�U*t���򸎞p�N<����Vuu�fUQ^p�*�*ײ�
E|�N�g̑m7��=V5pI� �b��������'t睳t�{NUcSJ=���,ڬ<�k�t�jh�Z5�T�1D �{��f�@�d�x�3�Y5ϛ7/�%����e25�1U0�!|��<G? �|G�	��s8߬����^�S$������O?z��7 VΟ�H�Ά����	�E�a(��÷�'���cJ��@g)��vT#XG8�e1�D@�|�^�z�i�:���	�Q�o�p젣��|�>��U�nҥSߩ�o�'w,]�U�\t��y�8U��as�	1�}4Ǉn��K� �d�KZ��Q���WB��E�X�����O=�mۓ��#Җ��f%�ٰ�'�!2��'���C�U<d�3w�4���js]	���fe������������q�iq���^�Y���+l�؀c�2�5��+�L��a����$%��b���d��锺J��nKSk�xd�@�`��~m����(��L�^��pq�����ý\�Ӷ�s�m���r;8F�U��z���ߵj9�[>�����o~���8L�����qoђ%�4����;�r�A5���h��{A�%�s�9^5oH���r�r-|l�r���f�ϸ��@���������G��YW�_o}�۔���Ɔa�r�y
q�3�	c�c ���A�^ۡ�����&�l�^��`K���ڮ��u|/�
�����*��s eL|o_�K#ĵ���e��|�I�jI�M��娘��R��j�.0�t��i�5���BZ�YPt֬�5�^�g;��m֖|g��� 3���`Ψ	�^-���S�W�Я�S5������'u��oՒ�k4y�U*{A�-ﳚ:�
u�ذ�V�N���e�탩>t��Ua�'L�Rʫ����o��)S���C�S����>����;5~�DQ��'_P6S�=&���B&,)��e0����j�ؗ?���x�k 2��:'�6f��zTŰ��ͦN������Lc&<w�����>$klX�c�$!jDG�Sź�y�j-w6��^P���ef�d�8Y�%����~I�Ҡ]�j5d�}|��ziɯuđc�����z�����+4c�u���ܮD�[��2�2����U�wr(cn_�ܡ{�	$����+ֿ�+���pJK����Y���i��>��Y�>������}�k?Ѩ�o�-~��;A������j� L6m}g�N�c����v�κ��{�|?��jb��cL�ܸM�f���͛w��g�mX�������
q��Aة�����}9�x��������{�Ś�O��������#ںu�f�:O7�0]�����3oԶ��pk�'LL�)�4~JgJa�!ޗow���^{��Y�A}D=]���V�w�O�M?O�B�~������K�])}�c���'ջ�H�B9��-��Y�9
�p�R�o� ��c9D�^��b��A�D�7�HV�fD������AQ;�ڏ�i�5ZK='����� �j�7��� �|�����UԦ�ل���ZY��=���}DUg�}�F�N���G+��t�����=�a�Tk)M�	O�4U����ne��yod0t���0^�|��?����jn���s�Ռ+�W�ԣj%�_ܨ_�b�Ǝ;A#F�JYJ�YU�4S`��r=.��)vְ����4����d���w�}�*w�-o��养ao�=� K�}l+��聾�0Q�'_X���_�����8�Q�G��jQ��ujj��UW\�amݒ	?�Z˾]���
5��-1�;T��OC��Ax��5Z������̪���1W.v��+��ھ���N��ܤ(�re�)�lP�R
;k�����p���S��?N�ʌ�k����o@�}��ڊ�	'2G$E��]Oe�A��(	��q����c���	B����T�յQ���RIjWt���]/<�^s�}Z�0�j�b b@�>�O��q��Z��S!�|H{(�Ϣ����Z�i��.��.�{�ijlH�ɫU2l���SU���^�;���K�P}#�L�Qq��6�U�>X <w���M&�;��S؄w&q@�^�r\_m�?8�b�����*�B�����+�iR:9J��Sc�p�j�&߽�iS��رG���C�O�@=m9�UkW�GV��!ky0�Imm%TV��h�v54���o?M�����&�"��ެ�z</!a����Ef�3G`t�6�[����&��:l_
�6�P��������c����'�DU�D2�B��5�kUw�08�F�*I��Y��H�bHN���X/6=d�ؗox���V�����];b��Ez��G�(ה�+9�J��	Gf\*Ѣ���&s�Z�[U��C"V!_	)�6E���PwQ�cn_DZ�c��L&��3g�����}Q{y���RQ�QwL����C<���ŀ��.��xa�I9lj��m�`�d�lZ_�(4Q��0��,���5hh�	Ke%�)M�6Kcǎ|� \���9b_�١{�{	�/[]�rc��Z���
ʦ��64��O�y�pr�a�XcsV�JU�JZ�dF���1~86�ٲ�������5@��s�̹aPA�^Em��ƞ�I�L2�L��</�&5TC� �ɐ�P��o�+�;x�I!s�d��x@~;��Kg�8l�b����f�~�xPU��������[�D8K��̏�C[7n���w����jZ�jc�u�$`U��-;c�<����b�	�\{���^�������*��C�Ր��!#JE�4�T-ըc�9Aox�[�/���w���Q�=��!i�#�N��3ژ�$V�)��u���%��9B��;l�����z�	�wY��Xs�1���Y�={��&MZ�'�m��	7���Q��>z@�vR�Г`��T�j�j��/�Ԙm
v(�BH��3��������s���:Β3�v�˲c����]?���7[-M�ri_���/&�eIԣ��uИѪ�s!d-�j�ꕝ��;U.7���3�1���)��פq�C�{2��ݟ$�w ���Z��Q%*y�SE���t�{�PKK*�(���`޺5����a'�R1���ȐmZS1wg�1��/~1��Lc�5���ט��Ǽ�{�����=�'��=�s^9������9(F��l^op  ��ٳg�8� <fÆ��ʹI�b.TQ��O�TT��U0ឞ|p�F��|�^.!I�����`r�9��zI��d��C���Y�X��ls���F]uլ���	����Z�ڇ�4rTZ��F�#_]Z����}D[�$U�5�k��ڛ�\��1�����O%�`fL��l�j�_����˦{t���5u��*;B��D�U�JV��m�-*����ԔN�����ZNJ��u�� ���BJR�<x�8��} n���w�뚓K�� �WٜK�`�Sٍ�c �[:ǳ�cP�R��R��x��M�8��=y�d��|����S�7M�6�m8Ԏ�]Y���*�dGӱ��%U��=q���t�P*�S�3f��k    IDAT�6iX�,y���Ջ\���Z���g͚����3`�����n��'���I��q�^wp��wvj�҂.��fuw��Zk
*�	��P:��VJ[ޓ7t��	�q�=�ϪV:�ؘ׽snԥ��T2Q��=�\������c4|䡡VwSӨ����H��|�+�O�	�1��l�%m����:+lr>XCUF���!���� (�&x.�p�����JYj��fJ��ZĤ_���a�fV�v�̘�+�J%�L>����4� <f���M��IM쬑/&�А���V5�4��'��N� �@~��0A�ri��v �E�@�)=���?��E,%8�=,���6wxGf3c�-���؛8b�QJ)ו�,{��t��g��NVk�0-[ܩ�fݦM��� \�ԩ�â�y�:d���+C��	�W�Y���>��6���{�����V�����>���UwwR���7:�ȉ�犪���S2I�r J`U��Ļ�Pj���
PdU�R��}�[21������� �ls��U`|�ƦL�(\�l����2����N�j�
?y����t��n�Y�	{�mG�oZ3���cgQʒ퍊ł�M�)��]��rZ�	S�޻�� W;�EP|:�DA�z�O>�d d�f��jh��m2�T��v���W^yE=@<�x��� kI�[���KK���Ԣ���7:���Ӣ�o��iׅz�;@xGQ�T�h�8�����K:wH���K�X�D�y���m5"������s�Yڶe���S����ZZ�wާ716�0cd��u�H�����  l����/�2�l�.��5��~0�x ��am�q~���N��g� �"�`��^���f�@�� ��`���7���~����^�ʃ>��Ae��m��7�t�H(IC�I��]��&�]�>G�-[��q�lH��C`T8�cMf�(l�6�c��^����4/�v�P��P��[��V�F���"Dvr�:ur�vI�`}fI�ۺ4w��Z��Eez������3V[�t��SU(4�"�	�{�	_��L8קþώo���=q���?J`o
��¼]0�a�6iԨ�n��Z]p��ܾ]w�u���!�����Ə���C��r����|T�/�~������3���g�s�'?�I��:ʁ�������^q-r�6N9��ٟ�Y���e˖ ���`��s��ζiv�`�
̨�<�LX�C�= �H$���'>q�����7to ��ܦbG^�v�ο��=f�^��"�Z����P2�A(�Lh�p1`�!��ݖ���ǵл���`� ��t����p����aՠe{CM6�+��<��CT�@ǖ-���}J���Ot��-z��������/,ѕ�nPG7 gBhM��p/��,�K����N�?E���m��u����Z�r�.�B ᖖ�f���f̸@=]ݺ�������:\7}�M:�4u�t+�a�	".=����6�\����
@���؟P@�`[2�U�\o�����??`&-�9:�@�U�#��3��6p�o~���S/�+'��'|��[���8?�u㉙lJM�-*l���<C���4����Z�z�:;��	@"0���y{Z�����#
+��1� .����f�N�%aI��,0i>f�ZL3g���,�ӯZP��Mw�}�zz6h����ʫ.R���z�՚:�usD�pR�DF��my�8%SDGTT��ل�h���x�D䭵c�ks;gm�w*�\d;6�Hj�kCk+W���gU
ݡ��=��W��|���o���-�'���l��#�Go�t���J�e��2��0vWp��N~��O"Q�!e�(+p
��7�b���WVӧ�v�N>��p� dmN�M�.���:̥�.~�r��`�t0�(���N��<o޼[�&<b������]ԝ�.�l�|���/~���\�� ��h��.�(<���Tl@����~W��կ�0m.0pp/<�쪊M����Z�e�8�aq��;k8��w^�d���o_�!�������MU�	�\֡)�?���&U�TQK�p�@��{��a�)6�;J��1�����"�����|ò��=��(�L�1�Z�?I� �l�r=���Ky��U���/{�e)QYL�w/lҢ7�u��S۰����Cj��ke%��Q'P�	������}V˄��{K��r=�~�<s�k��N�0hB�p�a�4�3�5p��
��/|�g�������o;���
sD*���}��w렂0!jlX�`��'�+EU�5�~̡�����m���_�,DX�,&L��g�5�uv	�H�8r��^�9���P}��![&	���/gZ��bc|l�Ahl���}��f�;c����9"��L����ש��M+�nׅB�E55�L�P;3J*�[O�7����ncfj�J;�vV����WVT|�跗S�����u�ܟ&�P[^��KC5�	ko��=KS���&Xn�r�mڶ������{�3�bK�L��(/W��W׀����0����-�?�;wn����W�vj'� e~c&��=���e�L�6-��f��0�AI���9��7�������L��G[X�s'�Kj�Z9�J}y�A�����ױ��-�Z��;Q3g^��|�b�k�7�~����+* ᥮�6tA�����da�x>R;� ��.�(�{�����6D� 8K^ ,!��$��}�{Ò;���	R�J�Q6-�z��mXV�|I+�n��om��S/e��׉�6u�ƍ=��9� ؄�|�q��+L7���)F�x����7d��p:�$���;���>]��i?���I�$$kZ�j�>:_���F���_���91���
#�+�ʹG�\���L�;bya���as&,��/�g��v�K.�$��(�M��ډ'���ް�x�A� T�;�j�S܇U;�8�29�����=�d�9�;_��v}f���D� |��'��ߣ��ڼu�J�r�	�����j�%9N?��p��A�'M�:Jx�w8����s��9�ӷC3���p�eP��=�RHX>x�/���� ����3�UWG��Ŝ��)<]P*1LK��UCK[HJ񌡨�� �
	��W˄��m6�2���"!N��>�]6Vf�S���
����r�I�^d����	>Ԗ�_�k���{X�BV�ZE�N����o�ӓ+��Cޠ�O����R��U�Pϐ��V�Ř����g�������k � I�*��m�g>��w��L�iچ)@uL���� m̞�1��8D$q˽��1��=��s۠�-�^��ݖ)����E]�����Z�zE0G ¼�����$��!cǍ3T��a�,3(t����2�����-\^�C����͂����aN�EQ/��H���PH$��A�Q�@TG�
�j��ɢ*�h�:Τ��I4�^��L�]~����'���z�:Q%����8+XA`
r.���1+����P�'	�A��%+^�#_���ڕĴPٮD�:UjUe����:b�jic�܆����)��T��ѕӜ��(+��0q�_}��!B��9��SO� �c�k��� p�;S�8c"�i�c��ۨ��<�Wp����q��3��
�ͪ�w��={�-�
�0�Q�V-l�&aFx?J�_>C�-��~���X��P@x�ĉ !a�Ȅ4�S��8?��9����`� ���Z�[Y#P/�]t�!qQq�Hl�@�uf\Q�RԢſז���I���H
xHM�����J� \Ӕ�3��Ã �������~����]B�V>V4f��ӡ�(7!���q��4����ڐ�Axպ���IU�傚�j��u'X�Y�L�&L���*���9�&\VR�>s ����ς��9⪫�
�"A�0����>�g�� <s\�0O=���Kd[3`��ò��y�
@�{::\���b�zI�O�}�݃�#7�\0J���{:��ԪCF����J��.���.؄q��@v��4��q{����YN����l%�&�%�� Ll<�=�%��
�հ���̆�X�����|n�~����ٱ-���
��4;,zi�jlł�!U7GL���^N+E��^�1'-O��񋱩Þ\;�,[�}���^ �d���V�3^S����l�X�f�}d��]R[S�ڇ�Ԑ�&��Ҫ�����>H�}�:�����@��WQ��	��:v��7懛o�9���8��l�Lw����50���
��|�+�r�����(!�S��p9n;4�`�&�����L�"�&�V�~�{�yP�	S�}����O���H�5F��ݺ��[B����%55�v��O%��a�6Nl,��=��H������;��܀V�		AЀ5�<0;��0d�H�6Q~c�L���jG�T
�Aw�>���*�rJe�J%�ܯW�{�B��I�T�M��d�: �y�;�#����8j3[�G3#?�o���f�^p�|lj�o��6d�(0;��"��0#��]���-�J���%����0bs�����Ǳ؁h��a�~|��!�����'c�o�e�p��WHV�nw�3���{�zEc�eD[�N$`~���s8�=��8}�m�A8��Ǟ�O�?/�}̠�7���dM+V���?�\G�=x����<]|񟅚�L�
��R�vmڜS��c�=��R�=�ݳì�L�����7����I�/D"Z��<���{�a���+��2� �I���	�x���L���yLÜ�aA8�o,��p:�~��{��Ƞ�1��Ft�_���v2���������N:F���i�˛T��sw�iϧ�;�&�'8��d b�AS�>Oh���_l�a �����*)q4��>8�x�Ax�ῨJu�F�H�o8D6����Y%z�5e�5�盂3���$l�퍨'����%�`�������	I�\�;u9xI'��~����'��<ϓ؃� ��������!;?׬����:l��\e�fE�wo�j��~��ab��z��������4էhl#7�������0�8��Jn�{B�
.vj���2�ǲ1X��v�ڔ��ξ��&������^���g��n��ݯ�]�A8����ݥ�l�M7O�ԩTQc�5dҊU�U(��N��(-u�&����=F�.�>�\sM`�8�*�[�2�����o�'Vӄ��^����&�6K �=��9��Y�C���>�{s�p*��ڽ��{Ӡ��ȭ�6�t���ܐ��O��:����i�Q�!��~�֯����^BG~tfANU�0�J�޿���&����� �����n#�'��3��L?!z ��z����|�T��%U��o���ƌi�{.<C�-���V,�Ԍ�7��3�J�Y� �鐬1n�X�ӕ`SN�2�k�>sG/H8���qW}�9^5�@h6䕀��`&�I�Ak��{�fñ��@36+<4?�7@���i{2h�1ӴYē�>���ǌ���d�x�?Ã����m��=��$���f� �^_���&O|'�� �qj��L�tr?ڱ���឴��oF��gE�1l`������"�?׫�6� �Y2�e+Vh��_P>ץ���u��v��J%kھ�����J=��M8���%�J7dU,u�S�EdU}{4�.ή�����#��E88
���г����c.��� �ؓ�+�>���w��x����&L;�+˲w�� �9s�|h�A�mÊ����I�R>�Ne'�	�x��B�U+VkѢ�B�bVeA����d<� )��x;��^f�)��{�qR�@h3#�|�|�p���\G��N�Ɋ��-�}�Mںm�.��}�P*����AS'_�Rq��զ�-'�5u��^.�F��pn%l�֎R@�xbz¡L�rI��X�<�e�cv��;E܊�l��f�?�gGGxBs-��خ��������0:�ȸ�eO ���cFƳc`5�5Hr//�<.��v���\�UV�0��0�Y&6�+��9�g3٘�ǀ��C�����y�N(B&1��qR�MQVj;Sd|O]��c��(�X	����7�Y+���.ї��E康����;��5����ݟ�>����6���;u�o�鰠.W�\K)Q��Q��`�a�q�	s����� D�^�+p��j�z�������I#��3���๏A�d�c��ް���|�+�1�|Md��j �{�w�AxĖ�G�J'���)jGx����z���j��	ڴiK��X�[��n�@a��	@�{l+[3{�mz�'OA��9္1Q<�< "�)N=��}���i��c�|�����sp���?������߭�{�3K��U����9������ՠ�U��kRO@�(^@�l�p�h�P�|>������sO��0P<)~����;6�&���`�b��1�`�2-	�=/���6��|h�%��Y%�4�q�������+f�1��;���.blvn6�d�-�U�Q۞m���� ����l�1�s�e+�X�Ǭ�J�כ��m{��?~���to�0�{i�b=����J�iB�c�.��L�x�+}����<\��>W�&�j-�r%/��Jg�D��)��i;~�O}�S�= {�>x@������n<_p�"#c��Am��q�U�My�����}�k}�����d20��	صaarۦ��!j՞��U����9g�+쬁p0�tҚ� ��a9F� F���G��أ� ��3L�a ��uυ��	�e��}ܽS&�H�Еל{n����<8�?q�N9��\�E�ϸ^]]��R�0�z����`U��8ᘭ�^�!����><�]��s��ؽ�I΋Ɔk扣�`�g![��#�0}˃ev��1��ywț��0 t*Ê�u=|-�=<�hǸ'�N��`r�ެrP4g<�Q{�N�dblfMi��oȄ���p<�|�mA���@l;d��o��(װra;|	y1��o@�,�y�6u��ܗ��/m�r���ݦ]�*l��6���KȌ�D_9��pQr���h�s���^5�AZ�)�	/]�D_y��ڼq�:�A��1K_r��nަ믿M�^ت<R��:��	jjlS��W-ݣb1��T�T�;�c�W���r3�3�hcҀ���`EO�\ܝ��=8�Y!#gV|�Ƶ�
�W�}������J�8��MSƠ}�8��6MjimJ��A=�l6�|�G�R^��mz�����x>�T��0����[�D��v
�U0�04��ٌ�k�[x+^��`�;�J����V-Z�s��-#���V�;�`-]�AS�_��δ*U��l�Y�t%d�%zkg�� ��b��&K&�MۘD '��53a\����X�Vf"�6@@��&#�8�}l�o�c�e@��� �k1<���J�����asO�E��,y�|��2�20�7?���L��9^�܋PĘ���'�0�xc��!��u��3q�iE;��ל�In`c�"s+2���Y�Z�f�~�����O����˸�Lm�9!� x  &;r����f���`O�#<�c��2`�{�����{�a��J�+���/�1mݼY�����g���g���C�7��S��TÆ�;�Oo{L�W�T�+�P�,YI�o�p��#���{�+f�?Bvf�V&��.�@lvd��EE5�-�I(`wG��G3o�s3�W��
3����aЙ0�a����*I�9loT��U͔�ΦT.��\*�
��&f��P��섁��!����N,x��`�R�����6U�.>3���F3�@��9o1ס��Y��˺⪋5��B��U��1�P��ZkP��P�rf�m9�
gP�>�cS/����D����xU1���ٖeM��FN0 �6@��D�0�,E �AD�p�m�n��&�FG���w�sv�= 	���� ���$���0(�e��;�0��m����?rR    IDAT� �.5�$@6�H�#�8����D��y�| 2���(@�〓MA�=��g,�8�������_d�,Q���x��w�Mڏ�b����}u�
�!}8��2Gބf��b��ܠD+�FI ��I3n�r��(e���嘕;�2xG�p1���|}��|ɲ���Ǿ������G?6C�/;7���������Rg������c���X�E�=�JT����:���y睁�!8"���0����u�Y�>�!3�nPzȜ1땵��e�x���/��(���J���;w��wܚ=��.�7"Dm�5ZK=')QM��= L	�r�j*��s��t���C�����W���IOL�����}�{�+
�Qs}MlɽA�>���x���0�W����t�k�J�lo���.�x�&L�d��&�t2!�=~�{�K��#a�01� L@��pfr1i�����a�ʀ�=��P���z@���I���	���c�� l6��� Y �s̑h���1 �`E�\�5v(a@�~�=?����o�&�p��$�� 5�gs��0`À KD����r$%� ��XI�=�N����
��K{9ӌ��� "
�����;mQ�\K���w��><��slR���{������	#o���j�%��! >���ڦ������ %B�b��W�����0��	�^�F=�9U��P��;��%�OWc6
�,}iS����o9N��c�N��L֓z�+��z�I �E��<�9�E���>��I�.�߻����~;�/$��܏�?��>�����tz���8�L������}�'+QM�)��� ��Hk3/�c��߱���	 <ӶI����&<Px�[��%)٥C�t������s�\�~��m*�S�8Κt�%S�Ru��;�^F�O�τ��g�2alo�\��Ť�@���yLT&�w ,��e��4|�? �hh� �0T 9�,�̓���n���И��;u}W��r��Afk<&L;�:�-}x +,f<@啓��PZV�6#01Q��s�o�t9x@(7�%���\�yȁ������� ������hh��=q3}����N����ʂsQ��$����F�|�c���W�[���{�3s���y���<�N��������Z�2��� "]�s�ua5�ɒ�ߣ��1��Z�f��ŴZ�G���$��)�TO�g�#Ko��1�)+��aj����x�m������[1 ��}����������9��`mM����- ��=��5�����@U�*=��ڤ�LM-�xZ7��Ѻ�=��޿UWGU�23�P�d��u���J&�}��uڶ�6j�E��<�}g�0������1�cخ�� Y���f�_& ��x���ȅ{���]Lfl���
R��"��59�`E�����1{uH�'6���)}`"��@�z��cF�@?m�� �d�� ��}z�8����N
Ϡ��"`�N� ��?�����x��ov~�^0_�L O�0p���C� 6ރK�"G���PJ���D����w���|'�ŃLQ�(&@�U�G���x������A��B��Y�)�}r�(VS<F�����A��3�/_@�1�R��w�:�4���Q����˵�2�[�U��������>���t�Wʴ�Ǥ�v���-�ܰ"�jثgcW��A>^M�'�ƠD"��x���{��?�=}x�������7�o|yA[���;c��t=: ���K�8|� eM��������G{���L���e��FtC�ح���GZ�jE �r�#T�K&��Ғujn�\��i*ժ�L�,LB�t���m�"G��
/ �2��ق�2Y��a��b�9
 `��Ra;aW�B~LP��L@�8�Cl�+���x �XI�T /�`�8�X"�	@�vp-  �rm��.�o�\ c p�]�`6�➀�}(���>� O��p-��<�L
�8�@�D! s�N����(-��= |��ʓ�Se�/rfL�f�N}��<���Q<�����E?�/Ǒ?�@��q�, �ǽ�@�PĘE����ȇ{�V�y()�j��1���x�L8U��W�s=�J����4���?�!�)�F56��ط���y} a�aja��w�.#[V�����$=�-�=���������|��0�o����W �9b@�p̄-�X(ql�;��`�'��.�53��¬���M�Z����,VO��`#.�XK�VmU2ݢd�Q=łҙ������:z^^R�+�/��b"���y�g��� jdò�A�#��a1�3a�,���d�������^v�"����y�,���4��1�Ñ6�7� ��`Ұl��؃]� F&|O;x>��P"+'� Z��A>�>0=;!�5�{1�A��N��L������	
��<��� ��1�hE�;�g�F��=�����M ��G~8�������v:���
�˸�Ǭ���V,���&���7a���٫f©������W��^SK�Q���U5f����c����C_�lC����+W��)rʦ�;~���66��fKc��{��,����8a[q�����nG����>���'��<ۥc.b�;a�	;��>Y�(�X��,�=i�@�Q��9��5[l�B�U����K�
�'S�+�)6m�-J(�|�T���C� �ђ�/M���T���d��H��l��fb���m�LjX8���o�0N�Cc�����M�q�	� ���
L`'4�&�X�k���8 N� R�t����㏶�0a��&;���P�PnY�6Y�{� p�M�<��w���:~����y> �G�0\��=`�0x�J�N>��c<����L �D��6�˱�$ Y E�B�M��6�/���N�y������$��߀=�����3pl"_��&.�g�=9�ӤdwsowLx��EZ��/�g[U�[ڔ�^�D"��l���V+��c�S&۬D�ݐɈ�nM�R�~
�a��g�8<�]�a ��@H����ڑL&�}���_�'g��5Llnp�t��}a�@�N[� c��Db��B���*�.���׆�W.�`�-R�M�>�LI��
�dB	�K/��	&*��Q�x ��0&'툵:@����6:6�D�c@�L�
83��d� u{G0��� �mj�m��^  �( � m����Y���B��m��eN;`��
����W#V�<`�9,�9F���=����8���;# �6���,w�#'�8������w`�7� � �ڶh34���_�k@���1����]�lA�]L'� xw��w�8oLP����L�h2�{s���=a�ƴ�-�w�wC_ c��M�3C�v혫i��z�G��Y
~��ڪa�KJJ��J%[՝��w�Kc��J-��
�j,��|h?�/+{���x��Zy��Y��g��a_o"��&�zd�Θ�>��^^�Z��it 3aw¬�,ƃ��owfwygߛ}9 ���Rʒ6��h_��Ɔ���-jmI����ư���Et�-��'�T��Q�]M�K/	f�x�v��ba�LL �� ��9*�la4�0,�kP,�c��!�����9:"L��ɲ���.C����� �a��	 A����j�e�Ov�q-��y�U����jh&ǵ�����h�8�u���9�	���̑��> {�Vڂ����v����z�'�B��.�ȹ��YA 3'��S��>��!|���Uy�p�'�w��5��
�}��(+l���A{h�c����Q&N�F1V��`�׮���#��\�*QN*�����/һ�}�ʤ���%57�M[�U��A�0�*0ߔ*�Bؙ�J��V�N$���V��_&>�3G0c�F�h�O�7q���}ʉ�����M8�>�Z+'H[����D^�t"�	aa�6w��Zd��A,6Q�K	w>v8q��߶+٫
��5kV_��_D����R:��a*W�����M�^�Ӫ���K$5u��!YO0[��j$�ι�3 s�D9�1���Q0#'� 8N&�3z8Ppvru(��ISbr��F������@�k�T�}�г�Ӗw��A�w�o�D����>�
��(�X����l�ٽ��x2�o+����J7^aœ<fJÞ��<1��m�W��4��� ��noq���w'�px�ɔ/["�Ւ��N͞}�f�|w����0L�B�::ڴ���̳��z�I�럶ܿm�M�(J��Ϗ�W�摝�~_~W1�M\�E�<_8���=�ұ�7[��7	QTs����W
$k$ʥ��eBD�!c{h��D��~��,�����w�b���$/ `qzk��⥃Y@�]{�}!j��j%�[����[��z����Mo�|��߽�^׾�c��ȆR�,���:uZ��T7��?;���+�y�Xi��/��������7��A.�,��c�B^^��)�tt ���q�Iag�.�R/+�|1 �n����w�;c.���o+���p�T�190��0�K,�e߳���e�6�N�1���_�|��+�݁���k���/H�����{�L͸�\%Sm�Э��vc�KG�=Q�v���X.)��(A��2���!��7��x|���v�ج�I��q��oכ���c"bR�Xi�!?�Ǧ3f�i�`\I�Rߜ7o�5Nػ-7�;��\����p�݉������f� �M1S�Ϗ'M�<��3 ���ۖc���`iG=a�t&�c����G>r�
�����t��h��az��՚5����ި��)M�2]G�K(����5Vvd�ē�6�Y�Ď�ͼ�8�.vDY~��Ks�-2`I����Vlv*�go�Ҳ-��F�d�f�?{g@П���Z���u���?>޷�U�p�~�ցd�������$ f�Ⱥ�.fx�] x�X�N�>��s��Қ�w����g+�N�����>�����ܷ��}�4�t�
ee���)��L��vY;��äͲ�j���z0�8z��m�G^�7����Y�Wp�o�m'�Y3�2�4t�p�o9p��έ��)���90�r��R��J��'qƘm;4par�`��U�i8`�q')xpƬ!��v,��h:�~�q�мf̘�g�'E ��T*���>���~���М�7���&jŲM�r�z�[T���� l��[+m�i��;�ENQ�ض�	�d���,������5��<�cVX0 �M�K���1V�����+v������x�����{P���3���{�t���9�+6������;�>0��uv��l�*=�p��][�>��;f_�K.9C������}���i��7�;�ao�r��a�M*�����r)v\�v�j�oV���@إO�`��ybY1�#�1��<��.��0��8̔k�)1�ơ7op3���ǎ�qՂ�bω�0�R�+J4�B����`� \Xv�� `zY@�܎�t�[&���2O"��]����G���Y.��eĪ��y����Թ�C��{���(� ������g��eK7�]��T�֮j��n��}L�� �΀�ϵ�����x��) ��o�a����l�f��2�HM��g'�#C�K=��\|����"�������s�q�������̹�;���|cv�/e�kNh�������ڦ��U�5{�.��Lm޴I7}�.=��f�s�n��^�w�2#���Xަ�Ɣ�lWQ�9�CD��x��ؔ��31�`�6�`���'59���qm�o\ɐ��T���
ګ�}
��^wۑ�����jI�".������	�1w��G�XK@�Ѩ�P���Ll�r�=���6Qx��tU��Fx�/����ĽB���#x��Ȅ�ӧ�4:��:+��f�}���K1�@}�ԡ��ŋ�k��7����0*(�p�c.TQ�];�\n����M{y����P.��?Nրh`�
��7����6���r]7!vJ�m[C�.�3���.fb��eg�����
��;s,�a�1��@�1���،gv��0�=y�@�����X�Ǿ�@=�4|XBw�}��N=G۶l�'?��?O�B���ןt�&w�����.���T�ϟ�9��V�g�uV�%|��I:�EH�&���*~�6]��
���́6IX������+�x�o
��p��/��?�V:�P̉>�m!:"W�Vsk��1N�&�4������fR#DK.'.�j� ��kw`���s���XQH�#�"�ŕ��������xІ	V+�\���wݬ\n�.�r����^���j��k�+`nQ�<u��7^rPB������`��c>�D�����˯���8^�}�c}_~�
������]:ۋmZ��$��企�lo�lw���-�8raW�tO��33���	{��}q�.A8Y��K5�#*�t�m�t��4m��x<�̏�K���ϫXn�M�Cc�zk��L$ECM�|��ɺc��6�c����o㋽�\�H!| 4c�ӟ�t�W����^�r.�?ĥ�L?��+Lp
�φ(��'��g3o9�5M"&���y���e/�W
'����\S��.��l�1�Mԉo����B3)�1 �d�1��7��v!t��Ht�����������,x��~z��E(������}:ċ���{lی ��u�?����z���*��V�\֦E]p����;kXKk��+u�Q�ao!}�^Lxg`3[�#l�I��[���(�3��Td{q��7��F9:���!�A�n��b�pVK����_A8fJ���f�x��&�3>�M��?�Y�'����p�utDM�V.����/��-�[o�����U[K�:�KZ�l����s:f�)�d����^B�j!�Q�^g#�	�NoBxΛ7/�ѯ��}�帆﮾��0���6[G�x�ސ-I=בI�8Nn�w?����0�܀2��duȜ���w�sO�{ｃ[�}��|��Mk���r`#J���:n�&O�4�5��z�kO\:n��@3]w�F���R�� D��sx	`
�E{}�������*0�_��^�Č���5aK�n�uޑl�7(ky5d����!�Ӷ�5�6�Ce��/m��_�B�AU�Bմ��M�RG�=��~��� ���۫ /�̈��_�r1+f���Px1�s�u.C�����D�_��#ݛ��}![O|�W�Ǡ:��&3Ƹύ��Y2߹nn�t�K��I�q����jǽ����@���Ym��HT�l�-\���;�jx[Vw�y�&O~��U|ERcS�:��Z���9٘!�t&2n�[��l9JYƊͅ�0E�w�y�}B*,w�����׾D�P����c�g�F���1�l�u}�wl� �7���T~��D��H$�Ycp���Gm^;����6��ՊԚn�ȑ#t����[�<\���9mܸ9h :e��
B�|BM��}���q�&�Ɖ��6��\�i�L.l������~��9T���k=>����=��Y+(��Ѷ��LKɜ2e5-_�]���W�6��%K�ӧ\�qc�V:�Pg�$lP�g'!j�����p��
�ūgG1m{���I��]��w���cQ����������TzE�?�0fz1 ǡ��x��α�|g��ګ%?�J!Ί����
�^��db�;�=sĪ%z싏*�ա�mM�|��:��w(�%�?���(�fK�����$�4U�i��0G�2��~�0'xS Lv0YL 8�#�3\��?��`^��	�ZVvA�ۤy�vx��5ϣĀ�R��3�J}u�w[�GoY7�9���D�sò���t����굫�Ң%!D�F0�A9f�Ih1j`�y�駃��n�Pb���g�}v�� S�?�q_	ź)�\��2�X    IDAT@9m&Y`;4z�ZT�ܭ~�_�e��P��L�j%�Jy�֯�R2դr��Z���UM�2K���t2[<�w�;[�ƀ�h�]��}����U�d�oX���۹����-�����@pꩦ�o�ݫ�	�fY��������
�����n���1��Nc6(�~|3�o�
����_Z�HO>�
�|�H8��U�ښU�w���g�E��S4z��T����O��a�k�U��W��v>[a�'<�|�M�b �܀�9+�&H��"Q��b�\l�3�����e��C&|Q����:��>��~ �<\�����}���!j�L�=�#�V�P����r��k+`�%ځAb�o6��/ɻ1���л��J`u�%xY�J�_=N0�jQ�D i@��E�=�b�SJ��[TcC��96m	EH�	v��	�w����
���O���`��'
�=�<���v�>|G�aL^A��v�mF�Ն�ӫ�����A�w��]k��� ��x0���!�mG�kT�p�!ż��n��l���۱+Ξ�#��Z������խ�tF5̉Y�6�R�*j�*V:^�)�*I�%=�L@���U�Ʌ�K��o��P��F�]�>�7laFr��3�-k0�)l��X��vk��W1��躐�ìA(�O>
C�,V�U@��s�νip7�����#7���R�>&�9��чh֬+�S����j����`�A�F4ڱu| �l�6��BC�N��`8��s�	ڎplϘ%0e0�|� �y���A�~~�ew��\T������B��v%��'WS&�Q!׬tf��h��.�eM�
c��1s��s�*��Tcd�l{��cgVe��5��U1��펾��ڸ7���L�;���<ۀ3_��ݫ}��n,�X�Y9%66),��8����O ���Ήw�v��/b������x���{��0s+V걅_R��G�DM��6e3 k��ʨ��j�����<\�dJ�f���3&j�@n.gi�1��v�m_(|�s,��{�E�k E�E&&0�|�6��{G>�]��^��^�3��Z����o}K�j}�@8�zjޜ�T&Nx��� al�8�ƿy����*=����_P��ҫ��p�1`�DZ�P�`ԟ5X8;/��'��h;�'�k��&����%�k�n��>�9�X��oK�͋E�|x�9�C0�Z5�bn�~��h˖5��ra��d�I�|��.ݢ$�Oq�%s�97}�e7�(��^		u����&>>��g�"J;]��Yml汼͢ݦxij��g]�j�h�nWv���y��f�՞cZ��#O Z��Vef��x�j���6  Kq���{��7�
Kwf�**fz�{�$o-_�Z_����uu*�(���M5�;aӃb1����\�g5�ua���sy0}_Q�|�P�����sa�l.K�m��"?�l�!�L���k�{0�T�՜�1�����J��^�rh��v�S�$��ٱZͤ�_���9��[�='��|�	�8�m�2e�~�_?Һ���UQ��8�H��e;q"6	`�A���Ʉ��B������ H�~�,� �ܹs������߅R�/����c�?���h��$s:`L��s�C!�l��_آ�n{@[6W��XJUKV4m��z��`JKb	�e��}���~�~�V`\g���o�|�X=�|����	���N�ݱս��1�}�l+�x%�@�(��\��8��e��M6Sp�:�*���}ضH�0s[��"���2�\}϶a�Ǹ�� c�s�&�zD�����]�)�]�A=���/{g�wU���]g�Lv�UYٷV�E4 	���
QDY�E����Z�B
T�.�V�\�hA\ؗ���$$�}���~�?�p�w&�dk�:וk2��_�y�s��~���tw���m�矡Y'q�`?�g��Ʃ����^R=[��|~�����L2��eW9��,ކ�x#&]�5!��"���� ��c����
pSmyĆ�棵LL���B���;{��%#S�j��$��h4���}W\�ы�����;c�m�۬Yvg{��P�lX���	'�E<|�֭_�j�2��V�a�µ_�:K�P@��\�a���p Z,�����ٳ����a�qx�OX8B(�]���ج��~��5( RR����T�s��պ�y�K��~����������k�<�0 <C�75����k̪���1b3d����1���f�1���m�ɏ���A؆(��l�l�F�G�4p,��F&8%Ly��d� Ą�p�Q�b`Hb�f��6��*� |��q�et���@��������>�a�8��%r�a{fɳ���w�&�e����B��z���n囊�h�:�2Z��/�`�U���Ԩ'��S��L�a�q_�Q�>餓��#E��z�	c+�Py;��
�L��0(�
��, ���W�}�,a�p��kO`��+W=��Q#&|͂�;찱;ވ>۬}a��Ca���3�x�	����*0a�#PBvj�v�Q"��'��}��G��k_��`�m������ �2�����;/�7HUÅ3���s/ ���q�W(���{nծ����9G�e\����^X%�z�T)OR����蜹��mӶ�1��%~5]�6�R3��و��04oAgl1�\��צB�N(�3��C�(��PF���CHG2�i���|�.�B� @�>3�a�� `�=6�iO�@��a#������
8����=ٸ�~���"��T^0�]s-[Ӳ��ۿ�j�&�gt��wi�i'h\���ݫ�>�L?��ot�NҤ�;)6����2�����Q~ I��:�������pe
HiE�+Ű���½������� n�̡d�_�	��˹�������g�;��5�S��V�\��]{��c^�rʺ�'�ˇQ;�z��춗�<�=��
����z�,�a�q-����\�b(
�b/`�-���=��&fl��k�b�$V�1(9+�>�Ɩ9v�`u�����2����e�]�re��~���я�7��=ۥYo;G��dU9�)+�9s� ᰅ.)쾙y�[���� oW�3kq��<q7�.�38b*.�v�7��"
rT<�_���/ڋ~9�;�}f���"�O� ?���7���'��nﲱ��6h�͌��f��\����������s��v@V\����3?��Q}��E�'�/�×�Ws�Y�J�~���u�u�V&;U�/�V�L�_Ŧ�����BzA�L�~D[b���7�����v�ϥ���'�0ǹ����d��0@�X�zꩃ�`�Ƚ�,��(e26�F2*�q�\�*����Ύ�Ps���c
�u��v��q��ÓڟE��v�駩yBQ���*��I#Q���q1�:��RlmF �hX�?��?�O~�q��!�j!t�q��^��,qA��dל'��]c�� �(uU�L^=�}��k��C?��{�����N;３��J��K��UTU�h� �ʑA�<���A�ƌ2�N���%�ڟX��1�C(7�I�7�.^C`�1a�1ۦM}?�^�H��}mⰾ��Ô�P�d��z�Ā�
�����L@L���sx©\�� .�|�O8�g�p|?���>�)�Pr�ʗ�铱yy
��%O�w���f�����|�9�M�бZ��S��7�S;l��.����^*3�5j*���U�JJ_���46��;��oX�SА�7}���?���&������:+�^3ރu���$���+�c<���8$��n��,�J&i��\������c�S֬^�V�=&�f�u��o����/�Z�R))������U`O,'Dc�}4;��VpPRL��ߞ��f)o~�C�0�0
������0�T؋�,:8���Á0���;�OިG��c�Ol�[.�|bX��~�zzra�rEQ.�}�W.07�Gl��ְ�?�{��� ��xO>@ȏ�c�Jf��b ���+ء�g]yW!F�%9}�=%��c��+K���Ϝ�����9�.p�qh&[�z�ސ�5�VZ�jc�}�Ke� 4���Oq1����\!���I�FhP���I�� ��h�%������jG\~�_�z�ŗ\��=��&N�S�_y�v�c/��P}��W�a`ja{3?1[��#�<*(y��ؿ�����%�I���<�`�@'g͚�@>L5�#��F�^��1�`A.���ųY�C��|�� �7�����pјo�s�k�.����������O�v�q��o�;�����Y/��X���
:�%Y�d+ ���"On�<���qز�\C���?�?Z�h� ��� R ���9w�DҮd�)��:_O?���͘��}��`=�||���=O��#� �`�3��HU�6w��O���X���8����钂C,`��Y�</�{�_�Ťe����=�ዑ�a�3#�k���LPқ�2��.3.o}u{��i<D��Bs���t�<�m֍�:���c�f�2 /����\��szn�
ݵx�*}���.]v�;����^����O�G�L��T]����w��P%��l4 /���,r�&�0?�H�͐7օ c�kƌ
��#���w�uW p��6b0W��3�fԮg3`�o"���cH �9������Y�p�c�S:�_���uDH�md�� 4���o9JG��Z�t�{� �X)�rc%�o[d�8�@���.=�oߏ�8��E9��(��Ua�U�e|�M7�ϓ�yIa��03a�>�eg�������J=����y����?+���V�\��k�aa�Nv1��9M�����#�ir�O�Y�Ȍ	c#135h�l֬8��oJq8�L��w���7��>���9�q7w�~t� l&N�!��Y�S�b`��@a����j�fo����6��9�#m�� �������)�I�ce��ιD/�[:C1᜖/[�;�r���^��Vt��gjC!��������SWW���˴�A�+�e��9� ��I55)���E��ǃ�K�/�����
� w�_���<x`�?���y�I���FF�����t��4�����>#���;���f�s�7^0s�̱ˎ &�Æ�wf6�=��OkK��e:٫v�NG�F��k���\��6���n����R�!�3tP�+�TK;��#�p���*��=��u�-����}H�'O8Y L&N�m�?��{�u�&��Q��)T�7i�ҪN�s��;�Tm��N[&;b��M�[�|%����o:Oxs'���u#�Y��8�O#���I�m�q�5f�CńcY86�g�0��O��z9�K��m����7֛8�����/�F�����\됆C^���q���G�����M`םv1 0p���} ��h�.��p�ւ��+V�+�~I�r���}��Ӗ�<VM�eut�����Z��_S��	S�U���,�ǩQφR�6.��4U��m��c�]j|�f��/�8x�dE�u {�Ћ�>{�t4v����"xl~�z�9k�!���b�.19��d�{��7�o�AxʚUw��&�-���}5��4k}�:��N:�-o���3��E�⣋�披EpD�)=Gp�!:��3�;wnȂ`Cq��|�ɧ�ӟ�tp�H�p+�I�r��0�es� ҡwh�6���ӻ\'e��W�ӏw��9�T&�٬Z&	\͙�A�{)�gQ�:���ູ�	�q{af�N���� h ��w�@g]2�3�t@����e6i����~�C#�g86S�-��Ôx�/~����Mq�3o��
d��q,�m�;��o0C~�g��]j>�����=\u���𙋔6%,�nݚQ�0�E�s�����+�>G�N;^��z����Fmmؘ��5%e���/��T��X�J99�֍�a�.eI���O|�t	9��w�������B����c����c�l��Ϙ�a���Y!�l쩠���F����r����d�)f���RO��CY6�N����k�����;�J��7T �Ӗ����i�v־�N�0��(尢�` �Ap�k����i#f�qY�$��u�[Hb�(6��=�"V���cΓ[�0O�֮c�KY�|M���6�j��N}��VwWC���ҬZ��Sg�����G<����H`�%��t��"�}��w!%��x;퉶��f��JG�'�}L,�cc���ص
,�F`K�{O�7^ȏ�]�!@ ���3���6
���33�o�_g
��.�E�c��$F{ i�0�z�F�s�{�k���X����>o
��b[��1̗ԁ�A�ٌ��|^���e�F(�_�k��x���d�IH!,�LP��I���V4i�����!��d���,+bۤ��xi3&�Z04ȋ�g���%F�c��� �C=4Md�z!�qhgz!_�1��p�����0�_,X�1a�&�_�#̄a� av�UJUm�������w���	a�Pv��k7�OO���"[�j�&�$��L���7�'��d��n��"A�ܩ_�Ǐ���uji&e�'1�f=����8�jU���ե9'�����;}�e�-�?���:-9"_� �d��;2f�G�v㝞�1���=:D�p�ͨ�<Zy�G&6��
&,��o�Hy,#/�!?��b��1Nڊ�a��nב���gB�v�����6�@�#��i�`����y�Á�#O=�yµZ��Ld} '�Kjd8ȳI��6���4~�P��y����F]��a2$�!�D(�Fǲ t٬;G�;r�%B�����i�����'�`E~ ��s������l.�8��
�x��ⅹL&�ʂ��p���f�	s�'�lM`�J�w��p�*I�C���� jf΄$��F�q��V��8�Y�cA{Ų�U�B%�Z�[��U.7)�oQ��S��B�Rk�z�f̜�l8i#Y���{F;����GNL�H��zB���8��8�h�06ncNXw�'���X�F�n�J�C��M`�Lf�D�5XY�&=�3ș�%�IL�Ek@� I��A�n{�6�a�� Mϓ��� �/`��C�m�	���%?�qzz��}�=�\ߡI��U+�(ñaY�T!\פ\�5��q:;�7̽z���0���f�p=��|@�= (�A&��K"��9|�3����f!#dF!3���⸱�o&< ��]s�5�9��~�m��#�c��<�1��Yi�K�"����PP*�:l�	%wƅ]���}V����|��SO����5���W_O.�P�\��+e劍~�s�Nꡪ�T8�O���0<n(#��$wZ��*��s=Gۯx>�	0������*�0ڶ�~����	�X����X��۸=��i�=�x���quH���L(�{7 Y8��3&�K0�a�a���c�����f@x�[Lyi~fٳ�����b�Z��U��J���y�T�*[��n;k���z�31�$�!��/��!/���CQ&�$���ymo	9y+�=a�4��������2r�VlD���=�=�rc��o��׭Y�^�=b8&#LO>[y�+�1���H�z>� ̖�.���0���v���K�A>V�F��J�[?�����g4���<M�d��_�bq��J5�
 <�Wف�ԯv���)!gLw�,�r�b��X����)�Ϫ?���c`L��~k�wS@�w,ް��q���F/�ŋ>gB��8��	n�Π����]_<�u�>�B&�P�<�������;�._�ܨ%�̼v�)6Ȏb�˟5�{zU����o���&�+����/���=�~���q� ��,�}��I=��2����EM�1����X.C��-�{�<��X/N�����j��L���P�1�k�\.��k���1e��׼����7��0[Io�$4 ���%3;���@���Yn<��3:O,Ѐ�������ꓢ�#�F���zC%��S�}D-���>E�>ݡ/����    IDATJ��y�W����5�a�����CHt�3����"p�PL��6�CyE[
�ai�	ב�t�K�c�����0D��`��&k�svv�x	��p��U�gx��Yxy>���x�;�`�}�'��X���W�?��7� ��8cǼ ������M��,��dɬs(���ҥ���۔���ڒ��Kޥc��3�l��H��/��Tn����q��T3�e[�� �/�^aQ�� ��`�l��cꐏA��3 �X;]��}޸C�A�`���M8r�ܿ]s�5�" �V�=�U��1�d�cR�Ó�V4IKv���`�.XZ�ce@x�u�Q@��;Pp��k; �"Ύx��������zVi��NRKKU}�u�x�����is/ToO�JՂ
MI���S�j���+��&�{^�1a�U��� @�:f]6�1��R����s�����>�$�[9V`<��3@ ��������	O ��kv�N��]XK������1R�.���j�T���g"//�J 0l��Y�">̵,���!���{��_B�rZ��y}�/*��Qss����<�:�8�8�F�e'��?��ϭS_9���I��,+�mW���z%�}�=x�v���]�*\����c��A<�D^�C�\���z/�ǀ�^�0y���^�ך<nc���l���]t�n۽����K ��J��Ϻ
���՗\[O�TS�x0cv�'pz���y��E̼�!\����f��ٹ'hF�u��O�-�f��:􈽴��U���:����vMF�ZS�X�f�</l��e9$���M��1 �S��
��-��0>��/v���r�7�o1�<����I����c�����h����z���AO`������ ���y&>�矋T1o � �k?��={y���e ��s aV���qX�g��1>���%�>�&�՞�e�� �r�*�~ۗT��W{[Y��;4��7�ؔQ��^������|Z�F��^��]�ϵ�\��X����~6����#[ד�m��蓳Bb05��`�޲u���!�� Ӎc��t��+
�ۮZyW{�/0a�3I�0��3�cf��'��	Sw�k<��'���v���oTQ3x�%�8C}]r�{��������U�/=' �SOn�;Ϟ���R.	�d�Y�}���"Ȏ0�e<6d�ԯK+��(��`4���c,��cθ�~@hF2�c7�^�3�T[2q��1��粓
0!�ҋ��V��d�� J��H����� ����Ʊy�c����r��llr�E���DV�1X��X�c�5^$%"a��8&�iC�ӳO-ӽwߩr�[���v�	�J�O���[�U������aG�H�}��vI!�I_8���k,��	Wz�ƞw�k���C#q8��3����r1�dan0�0L�l�\O�v����t�A��wbS f&�8��<ǩ&���	��H.���C�/�ȫћ��_��~��������w߽�rEI'�:G}�mR�5T|���'���f��ˊ��qrR�; ;����d'�V�t��bH�hDf�V��P 3b�,�|�&쉵5r�{	y���[�E�����D.�8}�3>�6���͡��A/$�� /y� �]rX4��&%�6�� p�(`� !lݛ�_5�L{�U2�rZ�r����ڰq�&���kߧSN>>��-�����2�膅�=����4��3�'dP4B�D� �Y�Fr,�'��=`���A�u ��M��rp�����.}磌�:oLO�skW��^�ga.�?c&�UR;!m=���غѱ8�.fR�	��|}�J������
<��0�E�;�Zx�U��#�W넒�|�Bx��z��:������)�[��S�N'�r�^7� ֆ2��D�)��L�?�{~6l�9�W�c���C�n�l ��Ӌ�2 |f#�1�.���a��O��X����������C����0;�`�;��da��o&?!<@�����=���;@����p�����l$!E�8mlH}dǨrz���oܫ��U�<��˯�K�4�Xm���/�F��2���?�j��?a�J�^U�%������4��Ĺ�c�A�n�����>�(�XZw�=��c]6��׫����1a�-OzaL�s/G�Y���Asw ��y�o
��~9��-��CV�pލ��x#?�e`]/�s]�n��Z=��O�������ߠ=��K��a��>����ʩ��4��P;��SN���,Ւ����WyQw��^�0X��D+}<�caP�X]���+q4C�#f��9O,_?�e���;E&L���a��S����v<�� U��,�x�Ӽ!�qd�7��4%�IZ&�)��8�J�:�@jZ�g+&!6O�>�\�l����E��|^�ƕt��h֬7���G7��	O���>���w����\PWOg�?C�B!�$���nCb�6q�o8=2�ݔ��a3/��ld��%��t��\�y�r��.\���1-e9����x��r�aÁ0�����]��c�A72�'��C����5�\�x��B���3�v�i/�	�n!1�Z���?z�j�U:�o�g��V�g�u�POOa �{>����C����B��"3�E!t<����d�Z������G��ً�+�|�p����Y�B�	�`FmX,����E���/�]�>��t�� ��<p��ɒ��]�B�qo�u���v�����'ǁ�qg5��|aT��w���s�m��oPss����b�|��d������?ޭ��Ї/�V�f�l�(4)�M�- L�i�6<V��i�I@�8{����vl�z�U̃o/\��}cz�F8����{u:V�'LL�ě5L�T3b3��:0T�'�n�y��<���B�e�|O��pD:&��S��>��oi��:�35uj��{���ɲ�<=b�N"��#V�'�3�z&��11f��&�P�nk@m$�{Dą�o'��<��f��'N.[���]b�.a��a����~r�d�m3�r��a@��7�:�d���=�F�v��]�)� 2� �yƄ#	��|��9D��C
��.yN��M�z��Œ���/u�)Ǉm���=��J=��J��4�����96rp"M���|���a�� �##�����66����8��a;�wa*/�zm���#�s�ܷ������9�~�u���!#�0����
��������B���=1���-O��@`B���cP6X�r�7����8;�q�
ɰR�Q�nפ�vjҋ�*��W[�6z���:�����ʐm��:��5t��yz��
��$=-)$���y,�x��A�1 !�ȴ���X��.��G����?ވ3�V۸C�gs�֦&?�u.�=�V�3�+�b�Q�7Ġ�^F�x����D_��ec
�dl���8LF�_�%|P.�n�;�q�pQ߂����K��2��@�*��زH�khժ����I�r�&L(꣗��S�E�:E�
ji��Ξ��[�J�FA�-����W1?Q�|�*��"���\wi|���3��u�{\�1��I���PQ���qaH�C$�W= �ߢ��A�����M��|��g��eԎ8� ��q5�#��~Ǡp�Ր^cpuz���t����W�bBL�=�0�p�����3�(ꌠ��Y�����7[4O9�A���a�TQ&ӭ^xF�dU�_�b�-Z�lI7��yuvV���T�t�����9� e-I�ګ���|c6ʢ'qa&w� ��cm� 	�2i0Ƹ�^�J�Gb�ǵ%�&�W���'�}<�@X�� �	@;Ǖ~`��k���o�8�.�@�g��u���ʞ!l���dC�>�o��!D|V��Yo�c#~�K!�Ax��%�p������>�zӛ�T�ҝę�ֲͪjm��b�8���a3T���ib�I�=�$�h��6'�5�c0�G6)��qp(Ƭ�G�a����wv�;��s�yޥ�N~q�ɍ��=�]a�!�J�,RԪ��fL����>v�hs\T3$ǁ�������Xx
�s=�q�|��'�|������S��T�{����˘�(G����xw��(mz2�uU+�����]}}T���">�RC�R�::9i�|�lO؜2w��|�5a��$�$[�_�?��qYD����4��e�͌f4rQ���opӃKY�
e#`#k�7�`$wכ,�61��G�"�!�`١�a!l��6sX;��l�� SH��������~y����Z:r���;�YI^�p���"}�Q6TQ[�b�����HU�!7�6�O�m_ԥF&�RoQ�ﰫf��&L����B�����dיK�z��c0b����7��x�	�S�X�d��xa�s�%�����H�Er��k��g�End��0�T@�Z`��{3coj����L&�\8�Lxƅ�m�v����(`^�6�s�zM�BU3^��������>!� �ԧ)�H�Bh6�Bz�:��@3�u��t>��yw�q��������PV~��o�&�0�c�9F���g^v�	�cZi�|��!$�У�>�Ro�����^M?I=]R�i�*UJ5�l_X��{�ٚ6m����X쓣�^�?6`���DQ`�;p���w��h�³�*�(�C"f��-�4@��|4��^ރ�xLlBo,|yK7zM��v`��d�9�� ��3���f `��9 �x<��x����`D�`ڃ�nX<�ט�,}��{:2�#�>�;ݭJ_�*�t��U����q�p|Q.7A�}d*�IS&�yCK�=�s�0�I�tE4�O��	�����a̚����� s��� �k��
+�'�`�]�ݞ��u��`$�4���K8 f,h+����˵�^{ј���,j/��p��b�®{����6�Ӳe+B���h�M�K�@�J"4�]g��5 ľ��m�Q�N8!��}�����gs��fፓ5p�-#�;��#f��3U�to���K����~�Ҫի7j¤mU�g9S$Z@x��P|>O�N�}u�178%(�A���j}�������|� �DcB�v4�Ǡ�c��Z��L�/nͻ�r��8%履�#�it]d���iz�d���M�H��C�`��9o� 0I�7��p����w�6��� �P>r�^.�X'�����%����kɲ't��U�mRS��\�W�ҋ��-�*�m����@esM��	ƫ^�"bF�}�P:Y�\�+��8:��@��tµ��r�[�s�}�7�ac���H,3��ZF�6�`��]�1K�����1�e�Y@��c��_�hۜ"��<N�jV��m:a�����{��?@ؕ��xfE^0�$!4�±���㸕'2�b���s���(�u�]����x�_+������ٸofo1��چ�*�6�_�s�:7vJ�����sEe�mz��U��[U�$i4� <}/��Ձ*jM��R&l�4�dl��3�2X�<�1ak@o�{̬�Έ�7���x�I@0���ۣn�;�>�X0�	�9�H��l	t�z�|a����:˖���?�i Y� �ș�p-2�~�=�;w�0�F�VM�
��f��UH/��?����5�vJ�JI;�8A-�R&�d0��8q;�|���m�}T�'������{�9R[ɰ���y1�~;���81���w������'�3�� ֐5� ����*{��g�l�����³����p�C��[�^��r�o.X��c�SV�^4%S �i��9c�~�5�Z�f��z�i��&�B�*!�3�!�V\��N��� �^���{Ă�"�&9K�$.��<�����o���ͼl�`�����o�)_�R6ӣ	��U-w�����{d�.��@�	��4��>��|~@yY�|��YO�f �ǘ$� ?('���΍�lDc��g��@G�0,���Ys��Ѿ{S���KX��3�&��	�sl֠�.X3���C��i���y �s\�g��\W��0b��;�U��)�#1��K��60�'�zT_���j��j*J�;O�f�\�B�v���ꮄ�����h��ev�����)��2����A��L��+d�gȒ�:�$ ���y>��@,���:gW�5��N��^̴�y>�s �{�'`��Q�V�����r�!��D�6��pso�A�����+�SN����_��~ul������r��s�(��M����(X���ٚ̝o�2���!��8���dG���e�	i_Ҷn)�N�nۢ���ɒ;ث���z��:y�{��פ��j �,���|.�W���dDff+�9ed�����-��a�5�y���5�d,y?���y�=*��h�vS�g�qYЁ�B�K��d3��j��/בֆ�9����@�(I��x�f�qxs0�����s�s�E>/p&��49�Zn��g2";��/Q�>M�ׂ�.Ҽ�OT��Rؚ[����auu���P�S����d�l O�s�v�X!/�
#�#p��=a�#�u�r�l����N
�x3�מxD��.��&����7^�䏐���Z�V���},�xLA��)/>������B1�r��ݷ�U�z�;�b�Z=���b�1~i1��Sh��`k'?v]qP*,44�ů��\���Ș �����Ზ��<I�܊��X� n�У�~����L�)sߢq���j�ji���U�o��j ab�a��K��pD±��@�UL>����B��N���l<]d�c�:���3y�R��}���� ���@!䙢��a������:�݇��aa��88�y.a<FdͶh{0~;B��q ����Hy�=���l���m>�b����/�V����u}貳5{����e���o~L<�f�8R�l���
;�Z!�̚
�E�O��zǜ�l,[���!�����!��v�w�y��w�yg��E1�1�d�<`������_��R�����{'��"]]�֢j�|���^���1�k�/������NJ=h�:�y���%O�t�#�0�!�Kh�]4&�Y�Wym� �\-r��c�y����F� /l��o��E��{b�P�L8��V�z�_=�kt�՗��g�N>�X]����5�G���y���E5��x0�/��9]Ӧ�|XGxɅ{��0�J�Γ�c��;��Ŵ�ٶdru�W��Qy�x�:���nh/`mjG�h�e�r�����β��i`�,�՘�S�(�ü��0�a8.i�-�0a�8���c���N:d�35�����d���Z|םa����U}�w�3���?y@��?j���.�kM�v��բ��%�^V6Ǯ��td������aLa���1�<�G�Kb�,ԓ����O�!ț�8)�5�9��)������Ż��l/�﹖�ID t��3ٺ_��j�|��kn������o���ֈ�5&�Z�hJ�q ��t�̃C8��?�ZK�?'��BH�0�
���;n��P����.��� ��[ɉ��x�A�l�@ ���g�pPZ��������p/��@���(p`x����_.�u�]���zXS��붯��^��nz��:�B�F�\K�u��9�����d�k>ʓ5�I`��} ���zP���Xm̈�DF{-�i��88�?�b<��{<�}�A�߱[�^�L�O�����[��v/��3& O�u�sp~�Cc|�gH�&�5`���x����yq=�0��L�|���-c/�� ��X�hb����V��oUϋ�0���^�N�|ʛ��]�5�������4i����G�����U.OvUF�ZU�BN�P'Y셩k�I����J������Z�#;X��?��p�����xA��~ثpx�ޅ�:��K���݌	�;2��}q���E��W]=L����~h�I�W�9��H�VUԎ8�0�t�,���/�n�ZUJ֓�5X,2|2�����ut
A9�������v�m�s^q�3 �-oyK h,��,>���0g���_�u��9vcE�qa�sl���S��c}�n��:=��o5~RC7�C:��Ѿ�q5    IDAT�uݚ5���4����Z�"'���	�MQshd(F2�Lw����l(��y�E]|��~;��+06��\��㉀m�B��G�V�5}��I�3�aY��x?� 8��6Z�M�v�g���.f�<P%��� ���qȇ��0ۀ�� �2�ŋ�[�+᧟Z��~�N�z7h�Ć.��,�tқ�am�.��=���~�}��_��4S��b}	0��/���<�f]���g��n�A.0�P��s�f, Ɛ1Ǔ�]���3�y��X��;�;9���	��������6!W�AX�b��֔����]~��z��m[�#֯�����P�Y�����ЬYoӯ��־�F}=����D��d�B�,OPB,�58l����ɂa��
�����{  ��Ib��(��t=a�3a/,�)�ro�nXx�~�˟��Cv�?|�Z�v�]�?,�9�H��Y5���
�e�� z@���F�1�RR�g��P�?i��f��<�q���s�ꭝd�N߁�X >c��ǘ�۬�qf���f&���K_gC��5{"�`e=�6
�k�x>���c��aWN��"`0��.�,�9�3�7�^�Mf��K�¥��\sD���"+��a�n��~���+��[յ�M����׼S�g�Ύ�n�����>���t�?�LW��)�Y�(�YQ!�{��Oh�e�¬R����w�;�l�r�3�����_���s`��#L�x6^��+��m����Q�QJ��"�E8��R�T-�͎=����ի�l+��R�QML�p��5K��G~7��!�����e�QB6g�BƲ $���_���+�8��ěY���e�vBA�4��+�NU�~��>�7k�LC}]���+�ѹLg��D��]�B�ӧ�\�s���[WW#ۢz-�l�%���
l	0��9�h���Ō��,�-�}a���e�¦fh�@����� l���^�ݢٟ�x8o�+��8�c�h����6Hq�G���{ ���g�5.$c��
=��X@c����3/�CΗ'���x�KtP�}{�<q���sk@���+���;Gtj|{EW]��r��[�������S;3�����}�6>I'$5�yT#S*I5$!T�_W:s�~�h3��
���"}�c҇�c�`��@5A�x+`?f�� /d�����H[�$Ƙ��?���z��"u�\u��fG����z�0����^����[&6���ab���7����<�(n�­ fC$.�LV%�w�:�zK"ʉb��0���IlwvĐ1�lM��F=��/��n�5c�.j���J���/��Yg\���&�5esy͞}�f�<0� �誨�Y�A��O6O���dw�w������k6N�b@J�S��H����i��h(�m�=�Ѽ�F����1� ��?��\�F�UG:/0D� �\m���p���w�AR���zb� p8A��G�M���#��Kw��ԳO讯.��\����L�r���e��k�~=��M�fg5�L
�*��Z��ve�lEO@�m��$-;"��q���n��"�	P�Ff�;l� 6�,R�LҐ��W��8��s#§n߃AMy8����1jGd��o\;�y�1qՊœ���j�Զ�zӛ�ӌ�����Jk_X�r9�c9E�Av�項���a��A�X*�j���b���ISC���$@���Q:3l�-�}��/+xb����j���V�.�L����׺��7��?��9���֯���mV��JnA�O>}�	'y�c�3u&���m�c �Cf�q��,4^�Ќ�6�k�׋v�o`6 ���e8��6�n_ړ�e:�$n}R?$�?cc7b��È!+Μ ~K|���`x '!�+@���6{�{��\�Y�?��p�b�̛0 �}�7�K!=��?[��.}*d'�<R̕t�U��ig�Z���T&�$�V�Xޡ	wUOO]�zN
e��jToY�<��x�7�����S"�����~7l%����L�!�a� T���K�"o��%�>1n�'�
,�X@�@��6n����������������ï������J=���1�L��M�Wo|�B��}B��	%g`mM��v\ǹx(�! ����ʧ+b�Z�LB
�\rIP0@څQ�Id��0�aet\��*�'z:~����R�Ӓ%���)�L��j�S���YU�7�����%G�$ LLx?e2ĞQ�х#b�f�]f�˓� ��.��l3�� �H��u�&�A������4 z�Gz�pߧ�f�N�73��P᝭iG����{b�3��x���a~3����N����u;���E&�8�Cx�� ��P�Dr��)����D���۾"��j�Kg�~��p�~�zT�R��MM�SU-OЄ	����������JT-l
���-s٘apDGX�!�@H��0^��g�&j�xӘ� ;��;����P�u#֙t+ި搩A���	<�ZO�����|.��k\;� �M��řkon)fX�ʔ� �qo=F�gLӒg��s�%q&�h,�`�B�3������2�ʈp�^\CHdF�
z��w�+��Au5,��7�blN%��`N��$���l�G~��֬^���^57eB"�fM���mR8����O �IQ��ד�)UN�3c
pܯ��-����l�l�=q�y�-\1�؜��k�kE����������h͜<C��t��c������
g1�m���/\�3`d>8������8v�wZVl�^���m?�c�2���z5iG���u\U�q���	z�Q'��}�s�������|�/�-�jo���W�#�X|���h����îC�+��G?�YT��a0���q��
u���i!��~�7 �aT���F.��Ƃ�_&<y��w6uo<&�Ԅ�i��l��O�*��]�b�։N؂��C[r�e,
�c(B'��vĖ�g��F ��=B5�5k��G���␄]A��1c�|*K��/�鬫Q�(�k���Y�WooWOR�2�d
�,��Ve0����&��هc��,��@y��o�'^��A(aČΟ{1y�/�,;������K �1�JV L�P����F `�O?�ϙ;��Pf�\k���/f[3�	��e�t�w�^Ω�H!��IA��6�z-��	���λ*_�T�q!Lx/��7��$Ԓ,&����|N��?��C���� C�ϟ���7�8���>��]���ο�R&cY����Nj ��󦒚��s�V�5�-_4���V,n���/d3l[v=�Z������POx��v�c>N���q,��1+�)����)1+����b���w�3�����Rc*y��6�%`pI�q�%��%1SE0��>�J?uA����
;x
M�/T	���Y��e4w�;4m�tr�Qݛ�~c�d�n]ş��nc���$�g�y"�8�~����������@<;�=5��F �����t��t{�S��g2\�m�G���� �t�R�v�"���.���p�Q���zN�B�z��!U���M���ڦJ��l�d�0�6'ٛ��x�,!�]���*��n;��a�=~0��y�w�DMa����xC�C����O�&^a�\�r �X�`�+�m� �dGP�'��ic�z�
Y�f���Î�34����+j! ӫ�\� (���z��ư30l� ��F�\�s���t��H�Â��f��_�������~WϯZ�lnɅ�Z�z�	�k��+��g4m�~*d�����3�<)=����%���qB[e�E�i�,��ʭ���{��i�|����x-ē��[k{w|�%�7Vc���U�v��QS�ګ�v,h�m�T������є)��cުw�C==���A�b����?��N��$d���u��s�v
X�6`^�3`6[�lp2��,�9�����kh�: l��^t�=�1u�w6uw�*jo�7z��ʚ2e�`]���mÎ	z�#P�2�Kl�;Wb��5a�7qa �;e��c��x1�v��n���r�AZY9c�^ߠb�������.��j�z������h��5��B���@8�����[2	�p�7�xW����t�3��dY���n��|�pO�������:	�^�	Cz!6}M����Gb�[�җ�
����������ޖ�{�{�f�~��>1C8Y�V�m4�IjK�I�ĳ�����m�x��/,@�M+�i�r��y�� ˜!��6b���g�p��3�#�Q<_�y6�\6��k�9މ������"�1?Y� ���yD���~Rq�"��gB5��`9X��2�@30�
O�1+-�5`L�^��B��Ya�X�W�z`�@�X(א��A�q��j��B�G--%m�C�
�%��_Tk�=�h�N�w��:��6� a�{���-�� ;�)F|n��q`/��13Jjz1�qrRr,� ?�	���o��1��� �e���L�8���[ߺ��4�|�Y}�+�%�|����/t�;NPw����W�>A�W�k�z��q�_X8�r��y�>��Ǝ9�c��U �f���F�����-��]�q�٤Ћn�1�@��;�I&;�:xŏ�׸�QL|��u�]7�g̑�6>"��5)[&h� �!}lZ(��8o��6Q�v�*fet� �n�]�C�>f̎�2�����ư�gN�I�A�����ߣ�v��c�?D�'��W��%%�q����*��� �p�ys�־�NW~+@��:�	����)1hDS~����7�12�j�1&�+��gZ���u�1�t����X&���Z��}�/�V*�������9��R�K�B�~��r���g5c�#��v{�^o��J�.��pZ)j<&�s&f�7h��Ldg�6�ۺm�p?P��8��Ƅ���B62��z0���]����F�]w�y? �㫥#�1;&Wj�c�=��8�<V�8��t&[*���3��}�N*O�6���1U�����S�A�v 뵒�}��Q_�����t�E�PlҳOm�ɧ�'��Y��Xb�[�^���:{[��e���Id���v_L3�X�̴=F���Gh����J��h�����C��بZO�γ��T�q���;��Wb���K�<���z���;5eJN�~�l�r�q*�K�����>v��Փ�G?z�f�<T�2R� 5�pO� �d�v����������Ƅ�ޞ�c5�r�5evmF�8�1�އÞ��S�����n�a���O�x~q{�/�0g���#��bU=9,�Vāp�q+F�:;ǒ� �w�xq΂��f oK���ټ�L�85 ��1~���V�ʽ������k��L�?|�cz�k_��˻4��w��/�Z8�4�rν�[.~iFb�ܰ1����w�(��!��x�c`��bO����Г�x��	$6��+1����Oa�e����x^��X�����4����X�z�]��٧���ޣ���v�5i��iμ��S�u�~B?���i��]4���{����2A��^g�_�<,5�qK�����):�T33]�nM@Lr�W/��egP������+^5��>�ûW�/��2��|�n���X�%sj���x���'�yaq[����ld�����+�����]c�Ke`J�Y��mS��O+v4������|f�EV�~q�>��k�裿R�(}��u��k��>���3T�4��9r��	N�7ڼ�5�@��̀��`�El�����ld����D����X��(9��]CV��Ɔ�-v�F!fk���EX?ӆ#V�4��;^��3#{Kq�ʆ����3���I��x��A�Y�����8�kƽ���i_3;��`{,c���X���G��sZ�d���vU�]�0��_v�N�}�:6v���\���
m��>��ŗ�W��-iܸ� �l�pQw�0;x��զ�U���Fh�~m���Id�\{%�����#BRvt�m�.�4�7wЇ��wY�Vΐ ��|����{��K^�G�_{﻽��Wk���ԓ���i���R? \�	�dan3JY����q�B�Vi��̛,T���꘻��1���d�=��1�1�z�!FݴR�3��Y|<��p���%6i#3��6ǋ7i���5����-�L�c�g�n����ux��������Põ'f���G[z����%��J����t���ּ�NPWW�>��O�ޯ=��^���ϿR{�}@8���4N� $AMn�W��u���A�����i����:�����%�S��M���'��^:�o8�jaœ4�vK���{�b���S̄c dW�po�.��|��kt�st��ǫPl����Yg_���A�>m&<��s� 3A�v�?n3���bOz����eo�@i���ǆi�g 6%��@�`�4;����wm,�GiZ/�&����u�q��:.���ٰ�š����H��c���4�r׻<"m�Y����f�Eǲ�Y��ѭ�W#ݗ�OCK�-��E�T�/������Ь�oP>W��zH���۵�#��|讀1�p�Q�?���4��$���s��z�`�n$|����0�Ɵ�=��0؀f���&��f��N�'�[��:9�Տ;�g�Q�qU�+aO������~��ϴ��4󀝕-t�l�������Q�:Y��,���ԱH���1� �l>�<.�9�k�� b��y���n=��o�(bvf٥�ᦔ5f�1�ĉ��i��������b&2T;�No�u��Y�~Y�}y="�$�%RiO��c٧��,6�d�I�e������D��!3����1��Z�sҞdl��bj[<��� �|ų����]Մ�y]qջ��YGhܸ�J��V���������M���z{)yYT6_V�ZQ��2�$�K_�� � l����H�X�{�P���5��_�翢 ���r��ń�pD�CVʴ0��ck���1����Daa��V�� \��Զ۶i�]�iC�RU���6^O=�^�x�ձ����/�0�-��>�p��@L|( 5Xx"yU��{贗X>�Ryp���'!���s��k�a?s�v��4��[����e���������:o����>�}�����C�q�؀�k�f�#M����^����Z>������>���Ǜ�x�J���,3��3����� �ٚ��x6�`�Y����>��$E-_(�T�	�w���=ڰ��9Wrr�1���#Y)S+)��6�H�9ֵ�H�H���M��Ga6kLY�zq[����@��t�l�(�$i �d�=#	j���<610��M�tJ�����U���d��Śr�>���[�yd�>��E�x�z��ԏhd5w��6mor��c��L�>�x�P�|S���p���"fαu
�Gb��.i���ń3��3hx �gg`����(1�1�4����)�!p��2`{\b6��}p8Ǚ9��a�5�vJ�A�v �Ά�����:�a挌Y�w���<֩��7��/�W��'�I΅���4i�8͝������Z�̙J�) oK�d��m�f�LQS���J���`��{ｃ�ͦ͞�B�)�wsI�����ޡ�<_w�u�t�Acw�\r�|z��FCeGp�=B�W���c�.���IY<!͔�(����Rw������a�������h�굡�i>WRSsQM-mZ�zcP�z��l]n�5wΙ�6}/re)�	dN_E-f/���7{��pb���}��J3]?�{CM�l}�(i��B�H(Ļ�x�����c���H�����H�7���oo5EnT�Q�:v7�vV���En0v ���N)C�.��i��R@�<Q��=���cEǸ�]����x`���Q����Cޜ�g\�ߴ��
��g�����/*��e�i����	7�b��PO���,5*�8��bSC��^�s�j�U-��:�����k�T���G��H�.��L(?��J���P�O�k��M�{S >�}t�s��B���	Xx�x���E����\6�"@t    IDAT �< .9�03-����SY�z��.yF]��SsSC}}��+W4q�d��Sn���
R�0�����~e�y L��2��� �!�%Č(�$b�|c@
h,���D�aƘ]��9f�~����� "��ras���K��ٟ�/n k�a!ŏ����8�m��|츞�r?p@���� %bx�Ϻݱ��?:D�U =�x�ϊNS��
8s���T���=��C������9I�q�Ɗ���U��<����̌�p��b8oh,w�g% �U�G�r_+��^ݠ��L�I[��TTSk���k5QV��ZhVo/ۍ��q�^�t8�ۃ1>>�}86����M��?��I�qɺ����@8��|���ߘ2a��<��([��B�0���I9A��A�cX
�,�5NQ<��}�׊D�< L^��{�A0����MM	&ŭb���[�1P��(�ٷީ���ڸ�O�Ţ
�R-�\�k\���ԝN��>���S�<R=a�>���A���4x[�.��Z�(iV�sm �ﲑ�Ԅ�a�Y�}1���s�x> F�*��� |�nP��ǹ_���:����� � ���\Y�y�S-p�sJR ���͐�5�w��FJa*ڈs�1l�g��ϸ����������h���Av(�� ������ (T�s"0流��G���m=�n��A3=��3!E����^eգr��9�/kVo_C��O�{�|s�j���M}�l�h�:�3#����/�)�<m���m`��L�^`���p�=2�Tb�|"	��=�^'��z��#�q���4PO���^{�؂���~h�Wߙ�XHKk�jՆ��ݣF��LN�����S�冝�1�E-BA��ꔫ�4%��A�if�Ii��I���B��̘1#��b ����G�v��@>_U�����[]{B�x�����>Y�>�<��7�I9�F1	GL�'�!&A�ˑ@0�2������l �FG�A)��Åtb�3[��5�$	�1�iv�{�:�|���L$�0��z�{ܟx�ĕ������R|�S�gr�����< 퀅`L0t�{�Q��Xo����C��<z	�@��u�6�S ��)�އz(lЁ���^@Ma�C�e��w�>���;E���.^�zU�����Q��K;m?NMM5��!&\�6i��u��ў�LW�RV�*e�.Ԝ
�$�P�` t/��2��#��b�9c@�c\���!��˸!_��(Rp=0�3���f�:��y�K�w#�����W_}��u��#�Lza٢���C�[���+�3�X����*j{�fO|�!m���Aa�f`e�H�d��Ը�>��;�4����5��E8������B���/|!���$�bya�@d��Z@�)_R��1�1ǙX�b5��<��]r�U��ͪJ��=X�=�1����ܟ� \��u�Pc����,���3��k��r�,>��y�G��	3�6�����0^�������� ,�8��(������\�������N1�0
�t�	0ia�0�ab9��w0�i���|Ǆg�>����y>���  @9 ���+���Q�T^�I��6��x �@tC»!����4�q�Y���[�C��p��O=�{�v�*}M�Ь�Ν�N<R���pe.ӦR�E����o_(��VON�A/���`��?��3/��<)g��7�9��c]5/��60Y�������1cl�27T=a��������{ǫ���l@���\sͅc
�3ϻt��/�\4�^9�R-)�ɫ�WSKKs �=�z��>������lM��lN�q>�7��(��Q� 1
- JO=arsY�Eh��T����[B�O������}3��,ۮ���T�8�+���o���M����i���R�@��Cج1�lM�w?�s0��A�ﵑ`���i �;� f��p^��ű������8��V�,�@76ʐ��bHc��Hߨhq��k]q���' $��K��γ�O�-z�'N��st�I�u���Ћ@��v�Oȋv�=��a��-�����29ai > ��_�@�0l�5,��q0��C���v���^r���0
��c�6Ң�Xo���z���s�"u��P{kNW]�>�=��z±�-�m��ڲ�{Z��YW&۬j� :l��K��.�{���M7�<��|�;�O<��`h���y��o�G���u�܏9�0n�/޸��r5�r<�x������"G�����n�馋��o��["�M֎ ��ٰzQ[����R���&���N����4Y�Oy���v=��s���,9�f}�a���Ą�pf��~����N�q,��p�
��<(?J}�y�k�UB�?�Ov,k�<x��y�Vؘ�e35U�6��?���ݮIo��Mݶ5���S�:�̋�ݕS�)�� ��i���*�bx1����
�X�Ǳ\�t�i��q
�9�Q^�H�2R8"�	�����@p&Ɵ~�)����7s�<��\ȡxU +z���5��	��q�y}���C(��`�.��;B��"��<���c��0�	`��:>G/��LpXυu����0fX/s���,��9j<��Ah�?!�{ˑ���� �乧�h�������Iͺ��s��YG����J����f�~q�㚶�Q�i��jd
�د����F������#dƸ^q���Qo�8�s�!��NcG� ���z��y�������8��$���{�a;�������Qq�8 ���~��7`LAxƅ�Mya�����'\)�B)���6���t��o�#�TO>�t��^f�h�]U��R� E�����s0��8��f�p.'fP�߼����x?����)[�8~�������Ї�SO�
�9�x}��sU(4�G�i�T)����0y��%������B�����p��V�����E0*�a�L���c�~�A�r�ӻ�Frg��c�n&LȀ��SB7ƞ� K�i�f�q̍�1	a,��3 {�9��yc ��|H� ����[�c��41���]E���B?�D�k�m������� x'c�w��ť��0n�H���n�ﳑz% vs��x>=��i�s�W��թ�m� �s��Je�~���u��Q�:Q��M:����y@�Y�������R�$��	��� )tQQ:� R�@B�Q�qG�QGfH�
�{g�5�;cEE�����S�~�o��9��rJN`֝�u���[���{?�����u����!G%�R��e���S��e�]�!8�b�40S�Pa���I�A��ڬ�3p}m����@�/�'�6�ߋ���q�8+�J9��>z�=�\7� <nժǫt,��nڬ�u-:����w�Y��z����ٙl�G͆��X�3o�#$�iӂ`~����b
6�Z�`��0ر�! ��1U𽽬�ۢ0p���U)���5���1=����k�F}�>�IS�虧������0�#*�L��-i��Q�'�[e�=�A���o@�
m0�s��km��@�s�n���¶����{2pa~ L�Ś�0��L �Qz}�*�E?-'�況P�3A�����Y�q�#��JPl��͎K<9ޡS.�ͽm��;~g��Y�@p/ƻ��k:r�c���B6��g�s�"��+���e ̭�������K�葇����ujn,k���u�Egk��պ��껏=���?X�}t��r�r� ?t	iJb�y�<�@_��W��6p�g١���?2¼ cb@���l����y7���#ք�X��i����X�ڛc�{�k9�N�:u���Y�|̠������?�е�X���">�g�q���6U?��h���P��0����a8��cDg�Y�`2��.x���E0<�C�0@�{X�:���zo��jG`��li���;tӍ�ʕ������go�[�v������U�U������9������Y7xt�A1��	���OWA��L�׈A86G����x�̭��`7Р�	�g�s,� 6MLV��@�Ƶ�m~q�P�ν���ڒ�	/�q&��;6�p?�1cԑ���dd3�ׄ����9���Q�C/�\�~9���v	 �N{��X��皱���s+C-�C��+��+_�??�U�^���h�7|Pg���ڸ~�n�y�~�����u��kn�aG�R�$�K-�F%�s�r����!?daYǋ-���6;X</��wh�<�gd�Yg�ٓE�9���>Y��+��3���g��= �i���	L8��<r��wlXA���u+LLW���� ��艺����Ц���7!D�d���6?X@�$ L��A�N��P�PW��>еM�	�c;jB���>X��dprj*��#�*��<h��C��RG��ϿI�-�������Kws��v�<�
��Qԝ���t��P%j{KY���0�OD&p���A�,�����bu���|��!е��&llN1��J��6�x������`WM
$9����`���C�T��Y��ǹ����E���W�C�`��_	g�K�����s�Ǝ�n�s�{���U��/�;���Ə?P��Z���jsg���Ň��(���15<���}�� �L/�>�&*k���b�.����p���P��oN��^`?��o`�&���D�Y.�[�VK�l��;��������l�w&:b�����sgiźez�O�14 t\�դ�	 �ax���N
�;2o̚=�	%���k�q���� fT�/���V��t��1gGV�a�WJ*tm֜[?�be��=�T}��3B&Вڃc� ��l����9"��3��cbS��3���O
��|��a`��8���06ؔW�X�1P6Ma�m��?@4`1��ǚi��_��@����w�cb��5�Ʀ����#��tQ��;��+�e�Wj��_W�k��[*�w���5�=*:���	����В%4�_k�}�W.�U��{�|�a��::��
���%�\4.�M�Ih�?��OA1`� D�s�	6\L���ڷA�"䎨�X3�0�e,d����R.���]w�qð��W�t��+��7Wߐs's�N;�T=���kɲ�!l��au�����@��`�ǃ@ '�pBx(؃Kj�4;c�Z=��c����q�Οv�i��.��%�os���-���ҟ�����cu�Q����|OIK_�Ѭs�VG���%�)͜y~a�\���µ c 4����w��?1Ǫ��A�ks/<Vsm�����LX���ju�{8���; �m��N�Ys/�^�G�5���s{�����ׂ�`�>>vG��ζ��8��h�zh��
ɦ�7�tipp74���Ӛ��z�wK��>G��q��ne�Ⱥ���T)�T*&Yq؄!bk^x�L!bD�xnجd�/�;�gy�[���0W��=�v�����0�
3' �{�89�lF���6�';1W��b6���Mw�����&L�ܸ�5��[�'c�舷�&�z������֮_�j�B�b	:wG��xP�^1G�[�����(���
��*��w�}a�
D���g�\/o�9"�x"�S%�/k:M���&˛5z�D���M������`�% L=a2��L��]�]���� �An�!FFqh�@��L��l��M��`�Vk�����^`��MO��$f�Cɥ�����5�m�����p?�9�K�J�ٶ]y���z�٧þp�Bݕ�s���Y�P���U�~��ܬ���^�ƾ.��\����A!�����&-��5���D��BRc��m�D�x<:[��v�����2�L ��	���1�W,���}cre�nظ��rJ��o�}��ӦM�8�P;b�K���g����<��t��g�W��^Z�2�1ǖ���A���#�!�=8Z�.���Y���r�uׅ����}�J��(�m���/�� ��@�-�m_�p�Gi��mzy���Ve2y54)0��Ͼ����_�ё؂�a�C'k���>fr��D� ������13u��P�C�p��X5�Y�ꟁq��
���MW����Ү��L*;bnٕm|-�m^�jY�Z*t��Tt�������fHDO�(��yO55�r�.)ϙ��A!���=}�����`�2����n"�K�1cF0;����{��̙�����:����;�@-��B�YͿy^r<� �p9��磏>����t���΄]E���9��դ5���4s����y=�̟Ö�v��c�p��!AN�Dh��@�`��}p���#,�3+S�Y�3��6�$��1 �U�]:SQ�5������6mH���*��qcv�K/��Z��v3��؄��>s�4�J�ⳳ�~zU��E���t�9��[˫?�i��sG 8�����֪ݖG-�0��YR�:_&�� �Kj��4�������l��*vwh���ҩN)UPW���B��1z�)gj̘�T�Шb1�J)q�Y�1�ݖ�3���μ�|@dy����GG�ܘC�B2'a�c5q �դ��O�+r>�&�{�������.��JB��j���w]���V�؄x�~:��)�(����R��x���6���z�bV���P�6G�9���{:Kܟc�<�b/?̖�!(�:�q��*�h�吨x2yңN��CJj9�wu�I�L�:�Ⱦk�a"��:w�y�<���A �)q�ݸw���1�:��H��;�m~qm�y��1���w��A#��Im;�N�u0������<�%��xQL���j,���ᯠ���W.��a�L�	���\���TW?N�BZ4I�'�|1qd��5&s��^s��z��fln�{�Ø�$1K� ���;���!a�1А�B}��_��0V1� -����&#'�6�J'�!j�̷�c�Ǐ<��u;����-���=E�6jB�	�a���o~��M��c@@x8� ?�,�4�,��:�<~#�{�w��� ���Q3D�I	�A��2��y��8�!���,:�&��B�[�<��
��rlwTج�&���kR���p5�J*���,��w��D���88� b��<f��q�c/���1�m/H�2P˯���}����<����As!��ׄ�ϵ��U�Ȅ������3=�yf�����`���x��C�U�$@K��|!�l�I�N��Ɔ&�����T	W��E�x,|mj8I֠��F�4,�^��l3Z���`8�v���a�0a��!m�9���F��m�Z8!�d��l.�J�\6��=��9���W���4�	7�7��Q�q��3��G+^Z�%/,U{{bǵJl�<�l5��WNm�{-�f5C����k�C���W_�C9��%��	� ݡ-�U���1�[l��Bq�~�����I��Sg��~C�ʩ�ҙ\���3�Sʒ*jea�I����L��sF$�jI��dj�X�g�v��;锖�\�i=���w�j��G+�KJS��U�u�m�}u�1o�GLS{GQ�JJ)�WJ��i��������R��K/�4�p�l�/�	��~!H�9��)���p�{�w(h���66�Ӭ�cC&t�����ߞ;w�u��c��qkV?4���V*�:d�)�������8I�M���Ͻ�ի��q �M ����0`�}̪��V�">���������b��
�*F!l4_��8;�͌�cε���*}:C���*�4zt�Ң�h�2���x���o�jU��� ���0�r��3�Wk��gD�!�W
�.Z�@ULu]~��q�)j�˨��H�Ѫ���^Q*3Fi�V��R%ӭ\:6�����Ct��E4�B�3gN��w�D�>�8߉~ ��sX  c�.�1_��`Ä��DJ���t��Cr�Y2f�6>B    IDAT&��];Y���R��调�����	Kt;k���!��}g���l�֭��}6^Yl�WV= ����P������v�|�PҎ)�1o޼p�PGTH{��߮�|�3!J"V�$f�-Ղ���L���l�F�ɨ��U��l&=��պ䒏�u;4�
��JF�g��)��1W�R�`����pL��k�H`WH����5�������h�u=�3�ÚuJA�,�њ�Z��G�R�Z�^�|-2�����K�Z�,;����>��`������ʃ=���������!`�kӣ͛�/����Ô�(�
^8�ӱ���W 8x��_�"�@�l`�Zeg�]»mX�P�uô�� 8i��V�iJ�I���ScƌN2�÷s���8�֋3&U{,3�_�g�(�DG �ޙ��B��te�`����C�j����L�ݖ7nX�_��:���:��7)�Mj��y�K���Zs��E�% ��1�P�	�����
d��&�W
����}�+�fRjn,覛/���:Y�9�TI뷿y^�<�J|�&N<P�JS�쳱�.D�
�`I�� # �@|�C�8̊��d�'����)TX�.	 g�9��q��sc �?������kሃ0�&*�Q�;�7�R�T`Ι3��ag�ׯ[Tױ��Α��-�C=�jW(�<��#t�'�% H�H-�l���#�P�����s�y�sQ#0�� ���:��x�� a��Pq@s�6��� �J��u�LݫB��>K�&�Ջ���}g~@�B�*���� 3f^��p�3�g�`^�WmF��hD;(�W
�+V,�c�������-��NU:UԿ������Y�^���O��1ǿ9�
W*�����F�f��0�ǹ;b��Թs熞�9����.�x����M� �DcqVᓊ��#ށ����)�@���E��.�qkW/_-�@�#BԚ٪VTH��DB�:��nq��,�S�(BA�t���PT��8�թ�t��2樂d�`�5]@���  �`&�ӏ���s6��hR�ahwΟ�g���&�у��}��[�?�R]xUH֠�O(����3߯)S�Y�M��F@xg����m$�J@���M�ڵ�ScG�t���k��wjs�z͞s�~�K�P��n��Nt�a�(�\}���d��#�a�c��Z�X���wp�S$����q�|r�q0���D(>;m[1����ua��;�Zda��*�e��4�8[N�ӏ͝;��ag�J�
�`��$麥LA��u���ӓlX�-gX�xKE`�-� /�W�w ��~��E�Q�ױz@�v�@¶'ՕԸ�w�������	g��ޭٷܨ^���������c�ЦMy����U.7�,*>�͜y��L9<DRT*���8i��H��p�@��RwG^������Ӧi�����Mw�W��V��s���a�&M>\)j:gɈM���٤�3�"E�Al64��.�|��7�u���8��q�`��7{�p�5Ny�k<�b�`Q����WųV�Ȱt:��.��7�[�n�xbsKc`��1WW�Ls�8��)D@.�B����u��Q�K:㒌��p�w�:�Շ��pC�\[4Ǻ+��&��j�^&�V9ߣٷ^��a��^���M:�Ѓ�l��:��K��7&�,��`��9+1G���4��3S��.x� ����z���RW;󮬹�]��3OQ�{���>}sѯ��}&��+����NRO1��!	_���͈�\a�q���\O��;v��������l��̆�̵��qDD���Ys<��,�h�kJD �zX�����V.j)t��ڹ���	��	������$����N���d������w�WBg��0O�	���3��.�|����k5��k��tj�y�ꃗ����F=��5��k��ѨR�Q)�Bh͌Y�4y2;�ĖOU4�W�17��C�8֫���7*����.��9fq�
�0��5TD�p��p�^�&Z��uX��q�'Em��c�]��>�~��,�=m����N����R�O���~���};�;`�y���qV����{�BZ�u[MB�w��0��'�Sr�!r��Mrh�N[7PL8�6����΂0��d�Z�`�J��ru]�u��������e=����_��^x�U�l��v���^�^9�;���/�����1i��L-���1N5�|l�O�����׋�.Z�ݖ������]�vQK���0��qN����������5�<p��W2l>0aq�m�����3��!��I����qi��vh��]�������Q�JS(>M�f̚��p�'��T+u���A�=q��n�\�Zu)��S��"��p��<�'iF�G�h�������l�LV�8�k�-�1=��Xc��xΈ��#���/0n?�f�p�'�.��@j������g��}�N���~�M�+m����<�6�ݬ*ŋ���ŋB�:�+Axي%!v�T(i�>y�L�q扪���֤��m֓O���_����J�:��C!����I����W��W��ߛT��oG@ئQ����\y��NL,�g��wo���+�u����X��'Z �>�@q�H��^f�NQ68 L��	q��y˽0it����=V�2��mVS�h-{�]g�y���f�������A��)+�)�*L���꓋ۛ�=F�q��/���;9�s=x���:��LĬ$vV8����w��^f���t𻁆�9�����r?��+m�6��?�q^L�P�=Z�4�\����̺�6G���g�jp��o�1�������Ƞͽ}_��>�{�c݋���0ǹ��e����scW��eID���.�4K��r�f��N54�U*d��쮍Kjo/�P��u!A#��͙�b���W��7_���gm<������ZY� cW̼��S�����+�9�U��|�Ec��'_��v_�jѨB�I1a�[8�zŝ��TK���|_���\fC��9�7��p|ߪz��vi�j�H�bSV�j^�BU+���K�/����*U3J��	�8W���5�����d��3�����d�i��'�A����,��!+&���kX����f��z�5�̽�Um���l��p��f}6�����m4�Ƌ���'&��^n69X}�/N����	䁺o3��������`��˱6�Y�f��a�bD�bY[�q����V�I�A�>�Mܖ�����#���bL�Au�4~L�.��]z�U�E�D�R��S}ݨ��y}]������f�&c�d,Jxq��3��qw�ׂv-��u��{o[�?��+vc�Hᜪ�	ׂp̸̰�[���9H�����ʃ�5h��vA ٢�c�~���Ժ5k(�r��r�z�*�S�ohQ)UV*]PEe�
�#�-���(��ʹ�K�<�'񍞔V�a� �����4�&����ӓ�L$��a�-j5׌ˏ��!k�~�y��<d0λ7��b�N�`�um�6�Ӷt����ك\�u���݋�˪���=��1+�6��5G�HUl��d��W;��3}����!O|�u1]��y�~�����k^di�Uk�(l��UL~�?��GWV-�hۨt�]�P;K�6n���{�Oz�v�c/e�.�N��t�Du�)�6���M��˹�������cR�������~@��y�Wu�Q/�H[���c�K[
�0�~A�6�n,>��b���U�xL��~haN�r����sO������IM���F�lV�RU��8�U@�"M����[� ��;k��h3��K�l��$�0Q)��>1	*�!A�	j(a7Ȉ8I�'��_(t�9 $��Z�����'� �qA���d�=U�l��b�]p�N��dbq0x�:��ɉ�Ǝ?ˀ�L~��K6��L{�;X�Z��j=�|Iq �+�^C��I�B;�XDlF�:�[& Km�h�F�i��XB&�.���m�t��yCO��g �\YA&X$y�ĭ"/�̟Y6ϖg��[�ߕ LQ��}�U�lST%^2!r�v��봹�K�:Y�l�r�d�qU*�{���	O��Z��s�x����rCͧ�߇2G��%[1h���]½���΂��
k üϷ����b��̭?&�C%�7[/�淿P��LU�Rw�l�ʤ���5&@�) <�d��a&7���%�� �~3��8��p���0)@��JR 79�8a|��\yw�1�9 ��K� �g�@1񩻊�)�xҖ_���xF�-���m���B �v�`��I��Oo[*Ϙ
ZLt�B�8��}�%�˽�~�\3��~�0� ����CF�G[��"O�I�*�����!��ܗPo��bĽ� M���:,X,T���; ̋E���vȀ?τk"K@��Bv$, /G}�4�+Ax��������J^jl�W�ܦ��M�$ �󅂪鴎<��e��ZM�.���WM5�.y�8d\ׂ�@�n{�����������= <��ˇ�9�Q�)&<��QadC��b����1� �؛��\�kS�j��?�C֭U�ܥ|E�[�M�ղe��kV����J �`���c�2Ø(v%� l�	 ;X�?�,3�aF|���9�&�yp<���
�	l  P� HS^�: nP@���H6��`��I�
�'���Yک���Ϲ ��u�v��~��<ٶy �̖{q-&�h3��Q�q�S�C�],, ��� <��*,<��s/��>Բ939�Ŏ�xN�'σg�,���^ 8l�c i�N_YHXmd�,���`[6�;���b��<{�gjA��^�M����c�}G�.JS�5����&�^T�浹s��~��z�[߭}�>T��U��3���9v�B��l���V���s{M��.B55��Z3���]f&Nx��+5�;O��φd�TgC&$k�����r���<B1(���*n��U:۴�X�G��"����L$۸��Ô��;?<��L�#�>w�)�U���ՓߨƦ������*��Z������Y��z0G�5�bM:�e2d�kA��2�`c�!�~� �l�]�:1��<��L~ؔ��Ӏ�1��<X[G��#�r<�@�8����y����� X�B#{���\� �xN��H�7���q.ㄾ��{����?m`���������S�9`gq��� +�8�|0K(�A.Ț�T�b���A���� �bd�����>g���g��u�xq��;��MH ?�ݶS�a!`Npm�X�I�,c��{7�\�bqp�mZߪ�v��}�l���ǩ���r�G�ι1ڼ9�je���VWwYM�Yu�t�:�����Q���Qf�|�]܋��X,s�`<ύC�)��e����������No�����4�|Otļy����/���ܴza}��̦Hs}5����P���Jp��q��OT�J��{6�L
ob���*��t�Վ������d@�v����������	�Þs�r�z��Z��S]t������^
;̚	���Fv�M� l0 &�6��H>��C��N�(X-�������W�@� ��f���0���G����C��^`ŨͰQ��8R���X8�@���� �˱�����xؓ�aV�7�����X!;=c �9�1ǀ H�1o�BΜ���&���ڮ%���{ ��XlXt�&�&�"�<Y� T�@�]a�L��&���dK�i}@saQ�"_�c¶g�"���ۆx��$ WՒ�/�-Rg[�Ǝ�j�͗�BX�t�ڻ�4n���v�mzmr��Z���U�b�++��w[6C��k��2 �w �,���f���LМ�#憝��a�&*�D�d��D���`G��J%��'|հ�0{��~���ζ��)�TQ��O1�W]CN�<�+%*��� ��#<Ջ��g�B7�5x۩��v�#`;U�jq��"�@�d��!?y�3n�~���j��M�[�:M'��`Vk�t�S�	��JՆ�w���5�� L�"|wu5;��	�2�=� A����dE^  �= fnL| &� 7&7�s`��x��+0cB0�`�� ���po�wHh�L��6/ �q�[�\a�,V�9���l_f�� Ф/����-Σ=��x�^��π0� g�q]Tz��
� ʹ�``�˸����3y.��p��EF�l����2d� [�s.L��3��3�9�;r䙳��o��bf*}�0h�:Ni��%z��_S�R���Ҝ9�駟�;�T����	=��K:d�������Ss�u�t(WGQ�d�O����5s5˷&l<�fc6���M��/�\kb��	��$yZ�&��e�}�	1G��r%��~��{����-�w_�baK���lu"@�R)+�n���'L�-�؀R�H�B�L�o��V{��v��F�� �J8�Sb�39 ہc/*�������)�Թy�����6o^���G���7d��S����_����JҖq(�% <� er�����Ң � Z��3Fd�V@��
�,lK�X�C^PX2e�H��°sO3E �g �ƦG� 610�l�@��!6Q �k���}��2 3�M�8�>9��`˽�D�%@� sM��Eơh��1���P��	�v���B;+���`��]@��J�3����"�2�9y�Ŏ6�Ok�Ȝ��\�5�d��	�̐?��5h� ���y^���?�+�l�KAx�KZ��UK�Jk��Ϳ\�{�z���ӟ�J�7��|OVW^s��8�DeӣT�H�2�T({03���GN��y�hO�ƳD�@V��ĵh<_�<�d��r��q<���D�geG'��:���W*�
Lx�A���n8d��Uǔ�Ǳ�Z!_
�,)��^h|��@M�vb�`GC�\<�a	�AD�a��n�4�z�:������78T�������N;P���f�m<n��ݺ������뀃���7�z���/�×~Lmm�p�Rզ^&|^ �lu
�}v~��&��ʢ�בpV�@�LP~�%�¶+d�JS�=�vu_�l��0��'��sڬ�c��)���ن�p��{  fl<&�:�~�xb0������ar�x�~ Q�f��G����1�Vo���N{i��/:|v�/�O{��H�s�#m������<g��$�����lwx�e�}�䲘�f�5�v����ыK�롅U,nV}]�����f�|�6ml�=wߧ�}�7�m�7�7ݮI�O�]=��R��d�Ą�{ĝv�i����(������a�4.>Ƹ����7� [s�Y�vf�c�@:x�g��&�q�K���{A��ٳgo)K@xb뺅�]m�3�\�	
y������+�q�����eU�����gM�`m04'��@C�`��j�đ�n���\F����g6��Y�A���C~%�|gE�n�E�?�+e�6����[O~��-[����a�{T��$LX͚u�&M:X�\W������=�j7�b�۔c�*�M0�����;	��������68��N�>������v73�Ë���+,3:O�x�q�l~�M��VK�����;'��teU���Y�q�9����30����m��2��W����Am �Z �Uf'����8b����8(�}6�N��6~w�`����#vx�c�˖�������o��	ҭ����N;I�m��9����T��{����M=�(�yerITQ�i�*j�02@���;�`*��8ϕ�Ȍ� ���������52��*�k��XC�q��@��,�D�`�w�5��s��t��a�Y㈫n:t�+d�[��A�!�uww��o�K���m����i���a(m�ST�Xږ��6ͣcѓ� � �O�l��7T9>�+_	v�3�8#�!��F������ǜ��+OG�    IDAT�+ ��ڭO}j���ԏ4i�x��wh����3O��%L���T�և*j��9��!�vN��.6G�m��N�X��@��6{d��r��"��;�œ��s�rA~�4l����s�����3�y&#���ʽ ,��g���|���Ά3�X��Ȃ����U_&�ߛM�U#{�9�?�JdO>�iƖ��N!�B�9����=�!��Ym�4r��zA�>������{YC�Y���SZ�b���Ejoۨ��Nͻ�]p�iڴa�>�/�_�ן�Ҳ����'t�qǆ"�
�d[#�Q�p�9��o���l�v�7�g��}.�5o��0v�����O�<L, ෾����*X���8��X���q�E8"�x���[���r&�}��9w��i�h�G�Z�`�JǱ�g�������t��S��w���Z&(����O���)�L�1���c�;�ٝY	��mo{[��~�{�9`G������������I�A�9��=�R��n�2�c��X�]v�>r�tuw�h��]p�uj�{[M�#f]lI$v�����Q�X�/��<t����'��fu� n���,/��|�sl*�y�A��s4��e�@����ф.d��	�1b0�������@;=�j�7�r���%���k�6��k��rl�����w�s����}N��5,��vm�#�ux�ŋ[��A:�%K^5���E�4�u�-�j�̓�M���_?�O��`�,��Oܦ�'��ik:$h�v�9���S5��1g:V�BB>>�<�����*����
��9�6f������9�@�߇gRL�e��t��;�뺩S�&����4m�L���������:{��Gu��}�;C��~��:;��
�xŬ�3 pf��`KF��>�h`��G��X_�@�%�53 �=�s-<�cV���chS�"���z�ձZ�<�kM:dM:l/��}�z������nVkkZ�*{�I���2:k�E�t(E�]E�]�� ���<�v>���F$�J ᪖�X����ʥ�V���C:�ijl��:�z��.=�41�j�}Qk[���L����جb>1���	���}����H,,���4l�̗���}�-� #�r���hD��W���	<6=،�Eڡh^^4@�4m|S�F'�(���J�J�\��;����
�؄'��]P��z<!j�i�6��N�!S������/�PHV�����%�ۅp<������?6�X��a' �����9�;Ǹ���5����إ����R�s����ܨr�S�GM�_�ިY��PwWV�j�7��f��v|��Z�gϬ��tF����.k��%z��QCz�T�М����oR]}^�tFݝK��W:�"�T�dT�P��v�b���0G`jt$��ؽ���`���7�	0��a��=*�^1{bv�s�5�X��и!�6E�u6h����������RK�l�����#�<rݎ�A�0 <�u͂����c��e�5�y�>��KTɕ�_��Ouw�H<��Vt�^fb���x1n�i�Y��P� gױ���TΪ��w�3���� #�4�#x��n˱3����nuu�V�ؖ�vR$k�U*JK�n�}�}]�6��	�>��532G`~�-�/T�1�����#Ǿ�0���/z����zM��%}����䓧�P���J���,��'�\Ɇ��L�M<��3qj�",�M{�ñ_�)�NҲ�Λ'{/��$�g��@�W��::�� q�|��l�	�����a&���OÄB���e�5o�m�s�1�w�Y	�c7�Z0��}<�ly����^�v�~�įU�%�/Q�a�?²��6A��*d����'}�8<�
v�����á�V'�Թ'������ Y�X��?�ca`Q�uVUPO~�~��k�3�UW�S6�l�Ġ��(�kR�C��I�U6�c;�R|;"x��@����;z��G$�+%`^��y-\�U�Mj۸I���'�|s���+956NдN�!�r%qВ�L)K�r�]3��π���K�%`i���Q4` ����7���XjL�\I�s�CS�l�4��\���8�,<�`|�;�	�'LX�\.�y�n�İ���+>y0��K=�I�8���u�Y�ӟ�{R/,Y6��� &:���!^]Tg� l������P; n:H��?:(������Fx\�$�jbo:�?Ɋ�.E=���*tC��J�;ܷГR:ۨR9�ԎH'�`�	;:"��� �����n���~WN��k�H`g$`~a�sZ�`�*��+$tmV�ԡ�F���PS���>5z|ؓ�2���$�48�z��8��sDQNl� N0�a�~�l'�v����û����\Nہ�>9d]:���o;|a���G`
\��.��A�j�C1��,�3��O+��<q͚���]Ӽ���'�E�z�;�ğ���V�8�L&�c_1�I�\���Kh���C�G��hv�qM �&ah�텈�`�#r�8�/��}�����"�=��p�t��?<�[{���,;T�kP�T�L�)ls��IBj�c.DG$�<Tt�P ;�<��ᶹbg&��9#ؕ�cn��e��N�K!���fحF��:��6�\M눩�(Wר�d߽�IB�P�$��[��Q�t�s��/��hѢ>��a^ޘ��8j₩�G@ؾ!;� r�����7�����IGP ��_Z�d���L�sn���7��M�g�w_�vas�sZ�H��ģ������Ǆ�e��T�0������E1�F�����>��!��f� 0�������#؏|�#�1�;�aV؎�f�i�P����@I�mՏ�oZ�f���;d����Z�d�2��O�	' |a(�CQ� �C8�2+�*�@LyWN��k�H`g$�5s˖�ᇿ�R�K�[�j｛�Ғ�w�[}C�
���<��������8V�=��	�h0G�Qi���cg��~O?��!��㏇�(�*k��8�YH�@(,�3;���9��	>0aGރ)�3�=��Ď�a�|���V������d�}���e�TQ������@xʁ�4s�=��Y=���}U�h(6a�ZbػR����Xe �L���0v!�;��L'�w5�Ky�)���i�Ɲ�e��1ʓ�̹q^TF+�6J�e2��K�K�����/��;�����*��E l��+��#������s^	��a�=�P��.ۭ+������ְMXH��ꐪSO���:5տN��(�kf�C�H�Z�`A o���>")�=d�X�D�M�x���;kҀ-�	�&�i!��%��q��tl
�0�����,�=��#jk߬2���.e�2߸��oVs�ԫ�?p��u���'x�Ͻ�碑.�0����~a.W�b���@��b�;��-dG*+a��=�	�� m�cUB(mm����Җ����%Y#횟}�R��Tvj���l�ޣT�Ki5���/��z��X	�V�	�9����\�{ߎ*j��)�0{�"�O��":��<�F��T�N��~5���=HF��e��B�j�G�M%͛w��>�uv�������+sZ��S��8U+cC��T��7"D-��>�����8I r�c@�;8�����N�ҹ�dġ����8���^1���3|��`@�&� �h.H!ף�z��.es�o�y���k� <f��Ec+�����!jg�}��;d=��ߪ��6��� �� �8V�^J��� ���@h�|�^P�9���w1j���"D����W��+ck\"*�#%,8�8��ؼR?����v�[�v�F�\�Z��[g��A�J�U�6&)�J' <�PeȘ�Q<c�ڀ�� a�;j}pL$���!x�}��#�-%08�Z�R_���*�ݡ���n�w�Σ�p����v���詧�뭚0� 廉��R�+��$Yc06�?~b��� + 's�'~v~,͊���7�9E�0����s�{z�?��ݗ�����	�v&&��`�����^?Tf
)'Y�;�nXA��5ƾ��|�	��LȘS?J�s���������z���a��}U�輙pl�v�\S����&8�!ܦ
۔O�&LX�� ��[�� �̜��Y`�0a�6�A8ؑTR.]��]�������f�#��
B�ٕ��>���T������i��I��5U	�4ү�����������Z�r�82A��#�	����/_JY�-Me͞�A͘�%�����|�a�ZӮ�o�SG���aB6��	c���K5 ���NlvJ��|���aV�h1?��o��0h�o��D��p{G��d�E�l�4a�9�{`��
6d�h�إ�z7	S;"��}���f_7u�Ø���ؽ}ݢ��'����F��رct�ߢ7|`��t���t�@���<w~c#ƏB� 1�%��x �f��}�C
�
��������?ݷ����4�v5���	��@�;���Oݡ�����ܻY_��{t��x�K������NtD�T��a��?t�z�����g�_Џ8�/�3���\t����xG bk�D�����t���K`0���׷���ݝ�R�-�߯3��6m�ܡy�>����/=������:h��*�K�P�.K텭���˂��5�*D�9~�m�з��H��Ox|�B�E�a�(�f��2�_�yET�\����a�r-k�f�0i���&RI�F�%[�Z���G��'��Z���~"L�8a�@���|ԡ:���	��+^�[��h��i>�����go�� 0�r��O�� $�>���"?8�"%� *@��j+�ج�.��,�RU��K��t��y�w;>�z೚z����3.V��S�ڒ�p�N3g\��SV6[��U*8�f��a(���vad�`r�~ ��ih���^Ԯt�.y�����70���Փ� ��Y}��o���U�ZJ�u�t�9����_�u�ݮ_����������?�9T�G���Nl�ٴ�����'l
��
iD*�O�_��onn�-���hB\a��m�Acv��_�4�'��wQ3��b��&,�u*~���e�ד�J]]��[o���iӦ��؄ǯ]M�Ɖ�	��a{�t�t����أ�Ӹq���p1�����?��`�&�a�AG1�s\�+k�1���3�LJYb��f�\�LV�/|�AE@�<Xo�Dz����(��on��j-_�gM�����7j���ֺu�:����z�e5�4��A�����c�)2��ׁ�6��4��]/���D_-�Woҍ�iD���F��|H����TԜy��Y�RG�f}�s���=�55�^�Ι�>$T#ĻB6]xU��}:0�ڍ>�1G=a���-���s�����:��#+�〯Am����C� ��]��%P���� s#đ�9�V>;�ӛ�Q����% <a��cʅ��ޜi�mη�yT��2U�7-��l����S8� V^�upN��f����F$k���7�G��T�{�VI��io�{1�ݖ�b�v�؄�֍��ݬ�z�N��מ��ԟV��SG{��j
�`�9+؄��\�u��N\�W�-R���"��1¶;8ݵ/���`y�H൓�� �l��zh�u�5fTJ��z�f�z�*�.��W�>���I���[u蔣�1M�1��d�^��0�
3�ܹsÜ_�j̀��������ĵ��i �d�;��8잏 ,ٿ /�؜	���L�0�g��qŕJ��9��[o�5Lx\�xb��
�d�D6�mN����1�����B�Pv�(�����xl2 0���#��@�]�B�	cv�m�qp��5�KF�6y`G��υ]<�쬑�1ݐ���_�{B���^G���:��m���s����؄{�VΜqn��H2�
�i+(��A�v�N�	�xG�D���+C���L#!j�4�Ϲ�PL�9-x�A廪7:�o�0�ՒVO��5�
��/��>��Ɩ�JSE��v��U%D-�Y�?f���p;s�p��͋`�
���?>�)��El� 7$�k��t��ǥ-}�XomD�wo���@8��>:w�܏�n�DG�ߴrQK��D�c�ʬZU�2�$[;1����!旕��sgX� \o(	Sv�84�������5RFWWO��^�u�{OOWXA�	'L;a���`�`�-w������Ru���K*�Z��6�;�*��4�PN+���sfhʔI��Q/�=�Q3�H��i*�8|��r/X�����Ȏ�F$��I�NHQY�V.	i�]my�4�u��W��oW:���fG������)��Q���Ja�V�$`�4����,X�Y�%m��k� 1��j���|M��/�7��p��zY�\�;��r��^����o��U�J���I5�;3�8�
��&Pώ����;4������ $�"na�ɞR�0��1���q�^޸B�\Y��V��W�I7h��n�}���^U�RU*KX]Uӧ�*���M���ԃ9���AB�9*����x�����H�l@y�5"��N�0�d����E��OiTSV^��t�a>aehl���T��Ln�R8�S9)ݓ��R��L�1�_ޜ��Wct��I�5�8�y�\�ak�6#�D%�b�͈��7YuXm|_��X�N�ӏ�~���+u����n�b�b�DG�Np��4�g�!W;��ǳw��ةeAqm����������?8��%������P��nP6EUa���F�Z�I�FOT�RV:���Q��;+=a4�8�@v�X�Y<�5�xa�ܯ�$���l	©���X�7*t��l����UU�Š92�w��u:餷j�}V�X�bU�$Ta�`g
"����-�y�0�dk4c��9�j��kƱ�����9��սE�|m�g۲ύ�V|=��L&��m��v�����k�*t�4Ä�ej�T�& 3e�h��r�7�c���ʎ-��8��1��Ât57/tX5SE)�YO?���=�P/���5�K���ZT�H%��Iv��sH[������PL�jmÎD��O~�`Ba��S�Qر�&(����#�m%08��li0!T�%5d�JU;���3� �f�l�0f�z�0�5�Tr|p�=sɅ����1�=c�͵ф�1H:2��ʿ�e��1q���s����L� �N��3����9�U;��M��|�'��}ͪE��0�#P'�
īIl����U��lA��@��<�=okU���!j0�r�]O=��
I��}�
9�ꛓ�wҝsd��8�����O+`LD^Yd��h�XW��f�#{��	��%˗�z�*���*aa�ʅ��Ad)�ޤ�R��@Ө�*���5%��{#h�	Ywwg�Y���f��&s	~$,�6_�q̌�ƌ>���p�&E�|��Zm>&�����;���W�)e���#���|��ի���X�A��qm���Z�N�	�(f۱m(�	W��ݪ����ڸ~�����rwO��+��P+�Q�J:ط���szm��Ʉ=` c��������Ӊ�F�v�,|�q�#��cF$0��&���p�C*vQĦS{���1Y�H��ԩ���1����G�=��W)5(��뫔X,���r98֞|2�Z�����kf��h3&i��c�5�Dc�#f��c��{̒{1m׀�k^Z�R�~�@�T5٢�/��f��+�k�c���%bVBǂ:���!(�f%�  �X�O�sN^]k5z�¾X��Ű��ŭ�m�_��U*��Jg�# <eʔ�6G�]��� Y���:f��w��,RC�p��	��e+_�׿�����7�NW^u����#�V�
Ŋƍ~��;	MjT*�$=�h<��|Ü�gBW�]'�I6>�1��6�������c��ٳA:h���0������y,���k�����Ͽ�Ug������W%pcP�����m�v� QO��X�<<v�&��M�`�<,?�-���J�.���~�(�_�\}�TNk�:w���`a    IDAT���G9�2I���ӧ' �#�����h?�7+��u
pf�%�G��q��w�z��N��A1�/�õ���0|W��Y���>�L�G.��ٙ�vN<v�����/y>���hVIs�\���y�r����FUK{hs[F�7�U(eB\=	��Y���5�xLHb�y%s=a�ۚ	�x{�qb�'� x��s�W~����&ĸ-q|�.aGG�*u��=氉'�l��|H�pt�qg��@v��$aN�p�Z�[���yW��5�2r��q�M%~o
Z˄����Ӫ���{�{���õ�����K+W�5}���jR��S�.'v9�ܙ�2irȶÑ��+MR��zW�����'C���svtt|�dlj��JaG��?�M�TiKIQ����n��ğ����{K_�)���[]��?�;�lyv5��kp�s�U�\|��������;�l���=nG�G������#�RW�f�]��[ޯ���%$cY����?��C&����N��:KeRɶ����Y��ɞn�i�1	ۙ>n��\�w��-��o�I���N�5�����keҙ�ϟ��2���5��d@�=�`K������x��44�w�"���3�p�2 �ٕ��X[��9�v����Z��Ԝ��iݚ?�sO�͟�Z��f=��Z�:�*ut7��\�t]6DI�7s��2E�
ay V@���ϔ���U]�>������|�eb�-R�L�d"ZM��[/r�N�-������F�����{0X��D�Ɇ��ҽ�1����}�xy ���緅�mӇ�a��`�����k8�$)+��|�2-Z�/��lӨ��n���{ީ*���G?����s��P�k>z��:�x��;�9�TnT]&�j%?(�������w��П�o;�I}���n���`���~o�mw_q�qSV�H�����τuk����0�R3a2� u$K$5|c;�iz���I��c�k�٫�s��wtv�Z�+N{�D�퍼l�
f��ک��\0Zw�y��9�h�^եw�~�z�-*T����<g��v�R�l0q*3�{Ad��3�-�[*��>��I�c hIo���m�3h��kGA�(�[��=F�w�~}�m �5���c���0�$S���{�!A8�pU����\m_���f�ܺ7����P18W�t�-\𠺻6ktKU���A���ܺQso����ȟ���[���iǩ��M�l&T%�M��Lp1�ZSA-�>>�d�� k?��$�^`̾��� ��cRi|�%�߻�ۮ�8a����q��Z&ӥ�M���۲WS|;�\/� ;�l��m=��' ^��p͆m��M���%��i�l,�t�N]m=����5a����懪m+W���PGw���z���^s��:[GN=J�䒌�
��w\��cOa�d�0ch���v�z:���Y�1���b��$}
��m���jp3��(ÔR���H���X�v���X�I�h�����HQ��=~{�E��ķ9H�v�r[�U���}���ѮQ�Ӻ��K5}��նi����&�ት:���u�e��ɓ�ΕU���r��j�8$��i7C���\r���;I��w�U����\�w̘Ì�EcsD6���=��s�a�6|�,�ݖc&L5@���\R��*���!�������pd�'*���+5x#(µ;#���|;WܞT�*�L����-�d˪��K�W����?Ձ�ї������?-�E�Fm�)U(:Bzr:2َ9�U��]ׅ��v�����`��̒Wt�P෽ ����''��&�W�����@̴������>��)���`~��]�Y�4i(�p,���� ��m�  �~�˖/��C]��4�Y�e�e:������������i��u�'g��#�R���i�V.���	T�2�؜8T;�s�:�#��c�F���Y&�h؄�Q�����xf0�S�{�����{�U�
�G^v�!�Z�,h��<��-a�N@8�K���[���!����aa�����l��ST&5�N� \���h�|^�öG�ap�a@!�`:�'e�舸T�A����wv���/WJ���+>r��Œ�����>���*����@u��}g���=^�<!4�`��5�9b�I�kn�[�q�$v�����@oi�P l�ؾ�a��Sj`�P�P���^����P6��Ȯ���؄��M@�H���՟\SJ)b�۽0DK�6�C�;��[����2GP[�[�\���657V4�+u�'+��~��g�������h��>v����T��Ov�	�l���0�0°�F��1�M�i͵�(f�: ��h�^��:��E0������7��7�����n�͙3��a-�~�U7�ۆ�{:�c��؄�J��l]F�[���Ïu:YU�0�Pi�0'������c����fwꩧ�z���8���/��{�e9��.�f�\��A�+�VL8SV�g��x�'�<y/u�!��˨�/k�ڂ���~�wfƣ�-�}�{���p�J=IȌm�M�!A2������w[�l���@x�I8�c���?`�j���qt�6����Ȃ��0���j�^-�m�{�/�dk��|3��(��o���n3~mӏ�@���y$�m�0����� z"��3�&�
;T,x��*���PԜ�.׌�*�+�����K��ǧ�h�����_�C4ԏR�@�U.�Sjm�1�����k�;���di�=䍲d����k��%a��l6���v�'�x��8�����${�Q�2�I?v�]s��퍦^��I�oZ�  �� �M� �����~�Lc�� �m*�6��@t��T�uvc����1w������c�=v��&�	so�f΀�%�\���U��Ù)J�M��{�Ǝ͉ݗq�Z�g�yI]x�:�R��T(R�>]o<����	�
��bZ}D��c��VL�wB�fǓ�f�m0�G0���1(hl��k~(��\�õj�G& 80VE��D�b�ۧ1���� ��18ԫv1��0��b^�z���_��ݪ�/��[.�y��b�S�,��ܢ��Ps�x
�r5��b��+µD��?�]�&��5YФ!��*8�\v҆�T�F4z��9��=�zꩾ�,��e���]
»mZ��9�y,NK�I�����3�l���z��a�"i���A�1x�#V����g��q�V/6�H���/���?�τ{�U	[ }�_[� ��N�@��1{7ͬ�w�*�jk_�Ɔ�TI
MW+9��x���o�ӓUUuJg�rw�6Y�nPkx�I�ϖW����n�֞X��)_
�℥;3)`xXM��JbL�H> �x�����g��6Ɩ��P&�>U�8��!V�X�ֲ��VD�1�}��'�%���,�Ύп��+~Nm�ĹB�կ
a�������F�]ñuu9
� �*�ej�x"��{�����I)��λ%� �O� �-�^��ܷ��\��I,ט�$~�$���t~0p��P��$���(̍�8���uu���~��}�qe�%K�����:���IS�0����j�(j���C�\����L�m�R*�jjjs��ȩ2N����\gW�g���ȁ0S�����TfK���Ȅ���P��Nv����ga'��  �`	c��M��p.�I��aA�e���q�]�L�:u�v[>��O��v̓�
��2�Q�(�?z�({�њv��Z�z�V�\h���=z�Z�^i���st�ݖ]�΃��`�l�	�bOfu��y��a~FV��7�����s�;6wl�eu���O��Z�v�Te�����ƌ�C�ֵ�R�*+5�Q=��{ϰ��{���ޤ���'O�؞h[ؾ��l)~@mY�aI:vb�J��!^�.I��e�"���8&nG�����&��+�)t�A�� �j�'wr�d`�a=\{7:L�c;�(��bU
q���`�b��$B���6�j�� Ό3#c��MS��'��"c�&�<b�N�p뢄����2�<qó`!������_�O|��8����6?,5f�-q���/*p/z�L�Ֆ
_�s��U��������=�+��6��o?�Xجa�(�D�ӄ��e���w��ή���Mx�Nz��zݞ�W&S�8��qT,�o	�����K�ro^0Q�a����wt����;� ��Ny�P"ֹ	���Ш�M ��/��!��x1��&X��6��'�%!ʢ��� ¹�G���k��'�]�`K�+0a�C���#���w���`����/���\~X `��:�4���J������}��U��a2�m��0-Pi��b���_���m��<�`Vm �-�R*t�d��*;C y]]�@����=U��/{�'gUvf�i[S6��:1�CH!�PU:�ˇ�AA �PE�E��B	5�Jo"Z�	���u�;��y�ݛ1����_���o7�3o����<�Γ\�e�!1	����Xc���J\�?���V��/�9�M�;G߳EwY)̼6�n�1�YW��ݯ�Ɯ'����8Oĉx�|l���1�
�LB��.��m
����A�o9��Ka�M-�7ӓ�GI�1aס���\���}�SW`��-"��.ס�Y]�J�	Yݫ|\��/.\ǒ�e�� $�]�u%qL�����qt��Ɉ;6@Ι����(�����g���Y�q���f�v������"�#�qEr�������ΊAXI	*r.����f���?s�!, �8�	�-�;�WX�p��o��Ƶ��Vj�7g�IsĀ�"8�����s�_~���٧���H���xI�^x��;��Q��Ր�9�9�?��!+��G�l�3*�E&f�E?��n�����OħL�p�p���[R��Ƅ���1��n�0l��x��iX0!2�\����ׁF��������:o���τe������K�������O-��|4��b��G�i�#� �͍`��)�x�|���4�2���cv��B�"K�@�A�<�aw���d�b�n��i�W(tXk���K;��%׽�Mhg��bN���9q1;���'&�	Xp�l���Ĵ���F��3y�v�r�#7Q��h����u�����x~�)����-��Il��t���p��Y�]���������M\~^��B!�O���g��j^��KznceׇRU<�����a5:�qH<����:	ܦ"�s�p�A`/vk��W��6k1o��;�2�x%A�[�S	�k������\_�by#����o!,��@R�Ϛ���	ekκ/��B�4��phqR��&K=�s��:�����&��_��5�y�d�Č]w�Ç7}VSY	���6,�B5���O�In�$���)S���^��)(�㱻ϟ8�Ǜm���e����[q���o�gќ[	�4��p5���H���^y�v5..�^����T�����e��鲛�c�=��6����(�����o��Ád9�	d�t�qqˣ�����R焍!��k����s�Q���B.��H��#W4d���>Y<G`󻓁v��0���um��i�S�Dt���a�d��N�E&78����Kf#UE�t��X
�{oQw00N)96L6K0��"�O�}3V�\�@�G)��~o9�c��e����<��F������T�0�D��ɘe��N������ۏ6�U�Ϧ❖Y��j�MQ�3�Pf���-�)�h�ùm�<�4U޳���˷��E��7�>�6T�"!�yw�&��O@��κ�g�I�):s��Yleˍ�)���E�`�M±�~�3am���ֱ���e	
�����,(ֆ\˳|�`�e��6Dm-�J�_Ѱ�b�b�$f�6LwL�i��~�3�u�Lc$�<���������_}�J�e�,�����7�4���0ٽF��׿�9�;��8��2�}Sfu��0��X�΋.��na����?����	��m[(9�{�9�s����"2!	�LI��JiBp7�JoaýѣG[�w�)�y�lxI� 566b�ԩ֝�裏ƨQ�p�W�.��ó��egJ�)?X���t��{�>�+�Φm�p��Yh��G��6cCe�![��P^�![be�N�pq�j Д�C��T�0�����C)ӈ�P(f�;{����,Í�kC $��������9b^�!$�Vf<��-����6c<C.H���]��.����\�%Ky��(����N��� eN��D�{<F�Dc�H;�sa���%���P@2�p�8S�MvW���L�������ܡQ4gn�����댚�Mn��p�?O&�+�ȟ��ʲ�9�'.ŀ�Y^?磫0��g�(_3�Y�,��ٹ2�Kõ�2�J�S�'����2i�*Y�Ry8IT"�d�o��ZfcXB,pL���'l}�Q��䇡��m��E,p#d����#95c�2�aS���8����ǒ���޸֙��O���� �,�ʉWd�>� ���_1bw\x��?�V�d�Esn#s�qm3|+|���������3?C�fe�Ձ�d�2�������"���3L�rPi^h�A�t�;�hM29�P���n�B���k�ΐF(���@g>v�<� \D<Z�[��B&�;�4f$@L��bY�$�vg���AT�[��}����t�71�yPd%0ǂ�1�x<06l�/:�� ��W�dO%�l�fs�NB1���f+e\�u;�N�عr�	XB.OO�[5�B�͓��e8qL�\+E˱�%45-� ��<i��5�g���NOfb�����j	dy�sx9&�{w&���
��W�{�F�nFZ�Ӳy�/c�9nv�n��5\:N��-��*��(9& Vŭ�T���?�.L�t:�{~����@'5e��x����:	�1B��M~_,��9G&����|5�<��:�1:ta��� �5(;�wY}���y}��f��,T"�CaB� S����'߷�%����*������q�Ɋ	��gZ��{y=�2���;v�������UЋ��t�I.�L!ي��嗝�X,�h�x��d���z�ͭ��X�.8��n�MN8s��f�V�n��9�6#�a����}�*(��wN�{��9�xѼ!���mg�曩|�4/��n��L -b~�i-�4��N8�{Ԇɐ�ߘ����tP�RϪe������3���O���մߢ9K�vʠ]r�h"�tXz�	:�r}�R������ �@eig�9&�r#��z�������O=b�$R�u�IUaIK��/�ʹl���mns s��4��A%9�ts��qV��%��>������ NĀ>=�@o��M�,Xf�6O+�w�f4�B��%�h��ȤsH�T[��6��Ǥ�Ǆ����K`�����-���X���bsk�ѷ_O��vC�݆C�*E�cP�ˆ�����ظ�D-r�<�j�1|Ӎ�e;�ܷ6�"�!�Gj0o^#>��3����������ݕv<òsѴ�(����·hk�!��6��Z{�(�l�"R��p��7��#H��fb�%��Pz0�76�p]�76�q���Yb�N�)��%����ȜĜیJ�x��У.�|��E��QJE�:�Ut��;g!>����q��O?9���4�ݳ\:��X+��ǐ);;��<�2ea�h<���� 5t�1D����&�u#�Aa�}Y̼:�H����B͗�9s(����H�د�l�N=��M]n��E����N��K~����9�x����;����"
� 2��s�>�[3�X;��ܹ���۷�>�n�b�Q;bܸ]��?^���s�	r�#�!P0v�7����Hy����,й���h��sg�Ճ�Nu�q���������>��c���ꪫ�5�嬑�T9�:��	Z4��	�?*8��꾻�d���i�jg�0S,�A"�g� g��x�5�$c�C47��F��d�+�УgZZr�b����_`��2�L ��{���N�.z��Ҵ��uJ�(|%�d�s5ҙ���V���_,���ev�5�<�$\�\1m��	^������e�����p%��    IDAT���"_�p���}p�٧b�&k"�ʡ� �L��Eʱ�b;jkz�����^�ioʹ��h<�w ;t�egS4�B���w��Ƣ���-x���n��6���@�^Q��D�Һ؜dEz�I��)�t�U���o{��L�Q��Uᢋ�ða�!�����i��"��"JQ�o'0{V+~��3��L]��^=�8��ð��۠��N>��_o�����Ǒ�U�W߄�S���O�9zc�q�ѧ���:���ɍ,�i��X���p�ݏ��߄L��G5���ß��}z�O�!�.搨�E&]v�E��T���᷿�f�Z���1c�G������kY��B9ϹYlPfr�	���^\���ٯM�M:�	´�����YSr�If�8��~{�,Ʉ�|�}�w:�h�I<���>��S�a�� Y����$#vQ�B"�|�9����v�'|����]4kR��y[�4�6�h8=����VA� �L՘i,t��yʓ*p$�e���	~���,(A�7��gJ�
���79�ػ馛:�׃�j~�Xa�:\���,Y��c��V%GÜ�T��gc��F��i�(z�^��۸&�b���j�z�q~�r*f�`A}���8��q⏾�d"�0��L	DB:G��������<Co�5��q�Uȴ-���7�o.;U�EDb$�=Ē`B�:��96���}�M�?�*,\�A�cР^��տ�F@UMK��B���%KZ,?�mB}�����y8�?�g� dM�h�?�;�\#�|����ȤCT��@1�As[�9G�~q�p��Amu�\6�r\���У��E��I�si�riԲWU)@6E����wN�E���b�^�S�������2��t���׺���6Ī��a��-8���֜4pC���y;b,��<��zd3�9]]M��B���5ho���s���}ɮ�6ဃ��ŗ�eV_U5=��҄H����$r�fD#Z�C���_q��? �gDK	��xn��r4� 
�PU� �#yh!�E�Q|2}~���a�Bnp���5�G��/\גDW ����1˰N�3�W�R�+�>�� y�G��Z%0r��QG6K�!A�~+̑�F�ʸ~�Ƈ~ءo���������=�S��;�c�Qq�a��*�-V]*���x|�ĉҭr�	�i�?�:�2B�䌎���:s��?�~�4a: x1��#;�7$�P�T�p8J���@�T��M�j���hq't!1α��\Dw8e�H?s������y1a1hm"b�_�u�)�����z�U#�m�5� ��C*�ܹ�0����޻�n=�[�a�u��̚��u���q�DZZf���cL��.�0�����O����ת�&Ç U�B6��g]�{��+°10z�!��Wg�GC�X���2M��1x���zۍЧo�m%<�ī8�UXҔC6���5{�ګ'bذ5-�z�&L�`f�^�D�
#Gm���kP,�ha��#|:�yV�����ӱ�ޛ��g�t�^|�~2˼�[l5n<��J/'�����Ȁ�m�&���r�� �x}0�0mm-Xc���醨�AP���;����X���q���a�-7B2Z�3fᓏga����Mb�m6Š����=�Y_���C��9!�R=�f��3�����BUUm�Ux���1�3����o���,"h�9g_��S���,��"|{�m���~�T��%L�����4�J	����t�:����}n�4��t��Ym�h����5�ć=���\�Ӧ���K��l3bK����|	�ޞ�SN9��f�h�p=$P��A��Hi�_g������qq�+.~%I�좋.2y��k�5ف�ε��q��g[� �F�>]I���d/2W9��Lc&�Z��������˟~b}�+�P�Z.�b�;'N�����?cH��_L�ɶo�L���܆�=�b�}��A��5.V��r�)���r @48�*��;$w$F;P��K��?C�7��.���p��Q�9?TG;��&�AO'�"�4�d�c1��d$��`.ǃ@8Z
Odp͟.�v#6A.�Ƶ�\�{�z�L�d�l�)�8�x^k >�t6�9�44-�6}-6���N��(~�Y��������-ns�o5��c��^���b�s~~��o�ek�JF��f�����ƚ���������Ghoˡ�z���18���Чa �|�e��G5hM�bР:\s��>|]�����<���hivyc����~�t:�c�>�L_�b���
??�T|��/���)�������K����V������{����������)�DX�>������Ä��_y#^}�V�y͵{c��vŉ'� I�r��8�j�Zcu=�����м�	����x�����j����Gs ��>��Gu*�|�A2Q�T<�?;2֢C�L~7�x7/\dRĺ�Ʃ���ѣ�`�b����	���=���~솸�Hā�>�<~w�x��/�0x@_��q�w�������I��o�F{:@�*�~��4�2�ѯ�f.���G<�̋h��|���Gu �Yo}����ޯ�����t�0�v��#1�n`	K^U/�}#q�V��KVvmq�Rz�߇�0�F��ɻ����DKZ�*�Đ!j<%	&������E-�Y�_�!�.C����'̰XFr1Ȁ�r�H�D���O�֌9���1��ɶ���,̇�S��2�v�c����{���a]���29� xC���!�exژ1c�ǝ�;o������3��Fq��%�s�YҒ�뮻����4Ox<�QҲ+͉;�9��K�Y��zEX�M����&g�:�z�1��`ܸ���k���������j�`޼�h�_��O9�}0�,n����%qsƤ��8��#�����s֯���o�&5������������~���/���Q��ZD#E��.~q�9�7�?.��j\����,�b��=
�����1��٧_'��$�-d���^����0|�zx������}�a1�"Wh�O�8�]c/?������tR�)E��s~�������<s�8ӢX�aqS|o~y�D��q�����?c�� V�&��[�E���e�^�{�~
�4��#�������?���C6ğ�<��ş�̉T]\�s0f�V����qٯ�-K���ޞF���<O��T~���p�yԉX8?�T�^�6�}�I8��=1�Ïq�����g��"��2��k��췿A�Ǚ?�S�>n�z��{l�_]:��/�◗�_0�)�$��x�6��.9l8�L�Ɵ�G�"5���֐�x��̂����p��+P�Ҫ`�q5=����}�݌����s0oN����lQ ԃɄ�E L��ײOθ�y��5��Ck��K/�O<a��.�đb
�$��R�rY����$1��u��� _r�wՖ �&>������z�vN�XG"�0��5q��S��7���k��7������t�Tס�.�_���k�=��:k�i���O]3���y�^Pi�t:q"����d�,ʜ ��3��w5������w_LFN0YCF�������{Ȝ<���X�I�U؂6�Jv&O�d���:�Pl��ڶ�����>���o��C�����h�^W^�'��һ����p�i��\��	S�~�s���`�� ل���;`7�g�~��r/Z��[�������x*�)S��鍨��l�� �G�� �=�������	�͘c�o��:��ʘ��t<����=�V,�U�؊ۭ�]v��By����x��O��=�z���N�ƛ����x�Ǒ�31$Rq̟7]��{wD�$}�9�v�ݦ�&SQ��iss�V���;�'����/2�Y�Яvt�>Xc�@���?pß���y�{��:}q�O�ƀ�x����g_B6�7Y��nɒ�a�15f4��<~y�o���_���Jओ����73g�#�����
�B(�h�B}�*���H$���C��ǟ2���6�}���/r�y�������OQW�a��l��y��X���6�c��������@x���8�'G0���0��� R� �@u7�F��ƌ���M�﫮�'�q9s�1���%��rK��rDe�D��EI %�u
�ZS$I���A�c+�%�����Ep$8��O��"�����~%FWP�,*��H��K�@[�K���~֡!�f�C�|�U$)�b��.���w;�?���\�H:�k�^���*K[�e��H�e0{�\�1�/e�H㵐�04�L���ed����l:?�L�p��Z���~�;�ŸH���5N3�������mI!+zМ.��K,D2JW�+&,JfN' �0Lۍ���ią�[ٌ��̌�\��<둘�a���;�Xlfu*�	'����ej.j-�!��X*ЊR��
�B�5ep�ͷڦ�H�=��[l����e�!��^��
%;�'�mv����cūo��X#Fl�q;�E]}5r�64�����X�Z8Ya�#H0�-���>�*��y�;dm~�Av_�7$��%�d,i�0�!�K�����0��|�-6Gz���~��dN��C1����JAU��Rֱ�\S�����c���a�=v��^
]]�\9�9�k�g��h�T5�z�I<��S(3Xw�5q���G]��7�7��_�A��L������,bL����%QW_�}���bNU�&)�N��u��IV�"��a��&���x���P]�n{C�1p��I�NQ�Gl���N�P�#_hCMm�eT>�̳x�o/x�i��ɣ���י�]}Wk_����(aE������H�3}G5UH���nSK4��G �c�ǣ��r��7�҄�Yeg2i��(7^j�����r�A)�H�}�9���[C�Ȅ�͙�F���ie3y$Kq˲bg��F��vێ�@tj'�%\��+Y�?�+Qb:!���ܝ�\`.vҥi���;��LX���|i���o?|�;߱z�<�@W�&���,'�o��{����|&�0M�]v�	#G���{�P���
�X���1�ic��.7�x�̥���ȣG�:��T;0M���Q���j-0v3Ӟş�x5�45�Yz�!�c�M6�D�D��ô�(�j{{K$��G�0�H�}�Nśo�D��a����hooEmM�|ȸk�YSRr������g�J��Ͼ���z޲��[-x-�r�������L�̤a�X�u�]k}�^=�C�ydŁ�ģU���N�!��1��af.d�����m�[>z�Hs~Qv1'pZ1�L���X2�x�������G�X$e���\3jj"V2'u�z��Z�03���]�[n�dCF�q�!Xk��(�]-�|ԅp�r!Xl(ɢ6��A[&�|���w��=��M7�L���8b�h�)茲�����H%��w�Y�)NX��-����kM-;��s���Zת)�26]���|�2�8~�R�E�$W�B�N}�׵�n%g���H�k��GC����s���;�k�3,�8Gi��^��p2����/>�[���c��Q*o��jy�ąQۍ��oiT��7u]� oȘF�d���E�I��aLa&x���f�>c��-�,���O3qȄ��T����yv�[�ʿWFX���06��λ����0[��w3�ъM�ooO{��2��wϾ8�cгW5r��9IYt�]��ɞdɽ�T��I����Cs���r46�d�����43��h9���&�4���g�ex����B�؆v�	;�ݫ��ێR��[X�n��W���W_�#�<jbk���q�Mb�vc�>�V�%��/:��y�����OV�&!%*��&A��2� ��;�[/&��z��������0v�]Q
�`� 7�(#,��Ӳ�-6�.���yx
�b묵6�8�H�V��4�H�<��}۞�Uch��'0g�b�1�n�e0D�����A�LCfZo�Y�ш���x�Ld`z4"hko�=�M����7��cϽ��[wT^3�>t���8w�RLRJ �i���?�g�}��	slx��#{f_�W���E�$�I�fh]�؈Պ\�s[�1���,�L�Y�$�>�E��A-�?q��@,�:��tApϹ���ne�C�?k�~?�T�ό^[�b,���ײ�gRv��0U<F ��M3Ώ�I�X�U;b%S��)b�0�$�i���IK�`� ���d�(myUO�/s|MM&��Qc��.��B����VኺS�'x�nU>x��0�d����w,�{�P�f��M��S�*���b,�l:���x5��̷B���{6�h0ق)��x3��ƺ\�6,PJ���x�W�۱�.���ݝ? ��5W��^JaWq�����w���GQ,�0x�z��P]Ͱ%��:pP��Jt^:	f�������Q��Q�C=ܬ)�"��X�,�+�t�v�w�]6�8�;�;v�
�@b��<�Fj��]�&^<��sx���a���z8p�Cѳ��B��`	",�hŜ�BM����1k�BL���z$r�Vt��/�"P���]��8u�b`R����<tޚ�������`�-G�gى,q�R�yj��t�C5)�z�	<�<#���)��V7��>h+���X�"C|8J�
  VY�hԞ�"0��S�	��Ĭ}�/�*�Q%r.�2�a�_B�y��R3!3�M2z��/��Ej��E���w1dW�fk����!���x�*�n��\Ԅ�g�6���;Ժr| �������k2'@ǈ#��.;u�׸�0k����\55�V;���>�t&�k�ջh����j���!�Rk��z�e�o�|7�)��X��s�!��Łi�g����E�$&e��5&����:�_�p \(�1v���N�:�-���5�\Y���_���NE.ߊ!��G�J]�BV�rV�c���X91~������N�Z� ��p��n�~J�r��e��E1���]�h)��v�;�0�
Њ0RD�M�D ,3EV���A{�ox��Q���zb�}@C��(�Pv ��v��Jr,�4{�|�1�.4��X����׊�S��2�T�t�rW���@ A�<x7�}w�""�b��lC+�K]�9S���u�ؼe�&"x����⋯�>z�,%s�r��^��u�g-'<׺�[��t�D�H)���"�:�i�������*0}]����~W�2Y�d¿��/~ԭrİ��f��ٓ��i2�@�@���m��紜�dҨ����	\��:�/O���f#���Xd{d����T�e�����oO8�L�%���"";ﴃ��O�r�٬�?�0�'�|��������'N:�x$R���E2�@&�C"Ve��`,w���D�=�o��g�GU���{ ��a)�"� �O�"�Z��=�-�*�?��|�D�El��6�c�q��zư�Te0�����xO<�(ҙfl��z����0�.�qԚ�������Ł�o�h֝���_�>���՚����u�ݹr�1L�4	���9'�����a���23�1�HH	B ��� %��ګx�ѧ,Ds���Ł��L� �M���+0�w�:{�,�:�6��6��G=�w?c`ٴ�$�"f�k5����x�-���{��p��6nl���	+��Jo&aD	�L�ȣTt�V9FO}��K&���bC���~��0֊�$U"\>;����h����ҤŬ�m����9߉1���o�r�y��K.���
~�g�{-�q�@�J�\� a %k�����H%hT�?`�@�Kf��KS������J��C�J�_��<Mؿ7j�����:��KC
������P��*�;�}�|���"��{��O�z,2�8k�DV�>�:چ%.>�����rf�j4)�a~Æu:)��Z�h	�@I�d�-�G{o���Uy1jv�aL�ȶ��:�߲�G]8���7^�3�<��v��z���}͂".]�[k�d�%���0=�}Ѣ���Y���F�:�k1E��[LK3"��P.IF]\��    IDATO�ܴi�%���{�յ(���61i���0.�*av���x���:���?�PTW�L
	�1�y�e.l"����3q뤛��i�1��?C�Ym-��y��PaW��Pb='�����R[U2eN�-�����:qƨc�ni���qh9�C�ԩ���^� a����X��^_���V������'>P�v�S$7?��O��O:�W8��|g�_U��Ap�������[�"+�Za��3&��c�Ǆ�@�L;�����r}g��8�J�
�����:��v$�I+9��c���ϛL���X;c�]�2	���+��և�&�5It����~�L��\CC_k�Ds�Be�.vR���R�|��b�	sF�>�N|1s�1�C:n���0z�XP���ddtƱ6��g����cx���p�[c�]wq H3Z=�:c��;�i�/��"�y�)��6a�����|wo����i�ńs�E	�w:��;&̤��o���fs��0x�Z��v́��`�\j�cA����`�;����v��Q��F�n�:�:4����x�W_S~�tu�Ї|� �ץ�%#N����Ps�����?~��{�/h�Ƞ���m���R��G�U�c�>Kf��1&v�=���!��[��-�ڼ����\��I,��4~
"�pK�>�����_�waiƄ��L�(�b�7 ���^O�����F��'�`�����U�
��b�>�乕����?��n�ދg2Dm c@��� l�˝'*w
޴
t�������BVV�~
�gU�A������u�T���d��׹x"Țcs��#)����@`�<g��aޙ��y띗��o�vۍDM�7�"�;��,یBgqmV$���v����|��6����0�5��$���='im�K$�� |{�[���f���κ�p����$A&�Yh�����:l�����&��ʭe�/F-8J� ��:�!�����|�m�PS�[l6���6p)WsN��~o;Ν�ޙf��'�����:��b���(Wi��R���@&��O>6g(+�54�[lf�4	�iv��|�"�ո���z���4�୷�FS���l�a�ӷ�1ב$�u]Fl�c�W��ioǻ��f��߃�\Á|YEp]��Ȯ�5#n����������ˌ�܃0�,"ʝ}	����}��+�o��6�Ë"�b�>�7������w���>+�\j��	&�ԭ �ى?ԫq��u��1%{���s-�����v���)Mƿ�=Q�j}^Y2~ڡ��ΤA��͔�8�?9:ƃ1�1.�"�S���5��+6�����bE}���L�B�ь�l�����v��&:�Lg�p(&-�>`�VTUV>,A�=SDUu�����QưMҊ)����k[ښ]�*5���3M\' 깱:�cîȓ
�3^����<��	�S�����0��=,�M)�oG,H!
6��Xl����խ���uD��@�E6�⅝%��*�=�v�p��+shl��64�%Y�k�i�a�."t�#y�-WQ~?�X��Y��=;�7Yk4��k�8vڣ����
�	�s9�9�)WX)� mmtF�.��"C�z���;V���Qu��#X�Y������8��J�}�O�ӷ�eY����O������ar6g+��D��Uµ�V
Fu�7����\{#G�+���+e���H��i��X��~�Y	��_���vl�C
�r^}�cuG����r�t�q�c��/��u�y��Gz���g:�4K;j��v�0����`�|�g�H	7�.j�	�e'�R���s���˭(���R��Ҟ;�
�w� P�K�"��pz�����d�K�#W��%���ʛC��7�-US�w1͝��ܚ�l�c[���p|e�	��u-]�}W1��h����z�����]!a
Q(r�3�2��QZ��}�\y߹���y�h4���	N�V&LM��a�X�av��!@��I#S]z�;k,}}�����^Y dE���Ү��U�B,��n�:�@��emB�{>�𿿬��i���X6w�������0�<�\|J���;�ry�]�.!�+3_*�ϲ�>�,Ӻ������蚻����o�g��i��@�oS}~��|�h���g�>��j|�N��RZ���τ�ͼ���:zy L�/\� �O>1_]���R�v�m���[�B�&O,�ں���\+�,|���	��]�ݲ��r2��}���X�;�騩�'��D�s��%�2��د��WW����_����9���|�>�?s��k<T���-P�wĈ�ch��y%�O�c���W�|�&|�y�حs��3o���6���4�r�����)��O o� ���=|�lK��nQ-�~�&�׽��YWLjy��
<W����8�;�oو�빗'��^�2?�u���l(��X�s�Y[%t5?���|C�,�T9����D�#T�M�$�h�?ʟG�/!�X�Y�ڴ?g���R��{�'u+3m��B�	��Z�</��k+5-$1�J�݊��R��`�;�����}C���et$��e��������|Y������q}r�U�Sy���돕�/�[lV?�?��_��+��O�8珈���	l�3�������
9��F��KN��R�,��s��I��֑�a�i%�w�7������.e�q��ޮ�F��Q�
C|����Vf��_���W�����W͕��(��sU]���"��b~0�@T���7���z��������r���խ��g�v�X��q��ܭ=�6��C�/�u{}�u��@�2�XN�P0�d`0�LqxLd��L�L�����Ϝ+M3��W5�W�����Y޽�*��e�mE��U�~oY�te����o�g�.��{�:��M�n�cޏb��STWm��L�+�%�7Wa�:)�H�2���,@ƚ�Y#|Sނ/i�|�b�H&|�E��[Ax��g�װ�Iu��m±�Ӏ���5�ʾ1/~��@i��a�(�]�|��T9〱�o�5e9pl����dG���T0^ނ�	�������u�/ouu��:��]]��t�	��*k��ݿ�wI�Xs�䎅���&��}֩a3O&�̤�^ͻxh?�B�	��|d!%f/�>_�G&P3��UӘ2�^s<��=զ�@x�E]��n�MN8s���f�R�k�jQq��V ��1�����f�a���V{�`�!��y&o�i��Q����,+Ț�
#Q;i�]u��]�۳Xw%V�g7��.��O�0������*�no�����#�F@&?;�����	�lgĵOF��cc�I��8C�&�BE�+,�E�`�`�5��B���bb�AbI<#N�K<�=U�����y ~�\�-�ܲ��<�֎��S7�;o�M=�V�PB*�B1��v�l�]w�Śpr� �U�y�BJxAܱH�Y��Ay��g��B��~rg#��L�gђ�>��w��3����*w)$�������J㑘��v�4��`����X=�� ��{��h�����@J�5u�T�u�YV�N���׋��'���'�"�Na{5Ue�3�?y�-{b� �?Or�k�q��*D��)&L�^v�i�4̟w#��D��
1�1z��ǖ�l�-�9VJY�m?|�]�D.��7�Ϋ�9�2�Ѹ�H�э�{�<�䯹�c���ؓ��m���G�?��J�p�k�M�_;uV�m�����-��.��<�1b�=����=(Y���+�4FK"'�� I�H�j����*J����ĺ�C��J��CI���5�᷑H$O>���O�V&��N:�i������0g=��F��9���z�V�a�м�	o����=�
��0�P?��7�B*d���s��hj3ou����47�ݔ�̎�,���&8���oM���P������zV���~H�Ȅ�;�<�)S���W^1��l�w4)����aGr��[}�X�/�j��v����e�[�8�7��|Q$�$�dƊ.� �A�}���� �gќ��m��Yky�]����i�ѧ���[vA*7I�+�W��5��;1ی����R5xj��A:��#�	Ҫ%L遍?�P�;�\~�pw�����3���#��� ʾ��%�p���Q�$��_�����2�
/��0t�P+JФ�K�!�v�������}=e�w(cЂg�]2r�����ly����� ܻq��#�m�b��Sb������Ǉ��?��#��7�~����y�d�܁�w�d���Ȇ))(�[�+�Ѥ'��l�i��&[%qP���Saq|�����X=��#�g���;�Зv�n�ă���o�%���('���M�GL혟q�Y�
;#vH��(W(m��S^��x6y�d�)|
�0���<��s���[/�2��Bǜi�o�/�o�Z��B	}k�X�چ<�ק�7w+^$���YQyi,�$��N�⋀��3�4�=��y;��q �w+��������d�qJ�)��|��� w���ek�gW����׎ q�k}�]v1ٓ��H���I��7#���0?O�ψ�A��Ad�����^)��O,cH-ϧ�3C�Ȉ� ��N�9A8�M�����#F,�2��%�il�!Ѷh/���N����/��q��oܕ(^��r�� i��	e��)�[�k#G�4`e0��;��q�g1}o<�!��t�I־��=w8�<�����`��Ϫߙ��Y6rU�q�qW���pHA=�@K�E�� ��{v��������"��ȓ-��s��̗���@�Cď�%&n����o�u���������ގ���b�L��s�9��
��ƃ�̽!ֲp;�`���c�=�������g��5O���]���y3r�|. �勃�}�-l� {�-����;������8h4'�B����կ~�O?��cpy����ᦩ�����.���R��Z�l�cA��ˮ30�Ė���x�ڳ�;5�/6h\�� �M���u�*��+CBW6qey��5O���^{YtgX+Ca�W���β�ӧ���B�����a�S��B+�@���
'�J��$~�	�%q��=d��AxqӒr��A4r���N�V9�q���ϻ�>�ގ!jl�2b�m��|���2>���fk����x#�q��͟8��f���r���;:2�)����8�ṣ��[����}_q��q����zt���0�l��;&��^w�H�QvSP1qW�[�r�B��Y/�Q �=%��`�)�篁/7�2�_��LE��s]o��&8ꨣ��&����QF�����]E��u�]�鐣����'Ű5ʜ���v��9AX	�Hi}�w&�͙7���,����Ϛx�O�n9���5�1קq&�5F�!��n��6�g���ן3&LM�J\�㖄A@U��&�@���]L@��ɠiV�'��� ��F�X`f�q0��@�m~���|2a�t�	�Ond�����pvt�X��B�t�DZ����Q	�r6̐����	��-���?wk�OY���������Ĉu�w�u@�r���&h0B���O�x�	�%��\�#\�N^-iʝq%�������!���Cak������9G����.�J�XL�x�ğvktkG�Y<떪�f���^d���18`L��m|:�S�J�1a^w��yy��&rGVlވ#�D�A����$�g��[o�մ���ƍC�^����<�b�<��/1�Ck3S.��q�h�%O��w��d�aW{�͌��	I���6���������_�{)�m97�^^%D}�+�j�U��/���c�=f�!��W�ċ�������R�$�aZ��I	hI iE�	����+�1;�x%�q��M�L���#A>�����v���3�l�s[�y�H��Hk��#�8����7_7&LV��߿Gș�U��w��F
B	��9m�4�9�q?��Qf޸^*�̸=?/��/��$`70}�~�{�i�1���v�i��[	�l]����>i�)�ɰ��Z����uG�g���(�9��Z]�]׷,�^�����ծ���8��LΤ5L��+��{�a�7-d:��������ә���/j�T�A�O�ϑ�1�B �02kFy1e�5��q-D���	�׽!j������ϟs{u{�1a֎�]��~�j����!Ӟ5�w,�0���
j�@J���\m$�=�`�.F���Xڎ��aFI��/A��#$�|P4T�G�+��Z2�=�uK��O������d3���b۩W�2;���_�u��d�����XU#  ����-"K˻>��I ��</�</#�ԉG;��~(�Y��zU�	�0�	Ԏ������<.�%��\"p$yLS�̡R��5�>f��~��b����h$:y���u+fg�>?�T�K�
#a� ��$��;`�m7Ō/>�������f7B�T��2R��<�
��	�a��<yS�y��J���Ȧ�"?�~�̕��#��PcE��j�	���;`e�x���.�l9��٥^�Ć	��Bgw[�-Hf;�կ�#�*G@ �*������Yl�Iv�'d�
����U��N�{�)��}衇h�5~v�t\�W>(���+�e��~��_��&��A\2"���0U�̚�wx<5%�����ǟڭ �s��̺���UB1(��1d�:�k�=PSW������wA`���0��@%�̙!&|��ݎ@;v�X{���u��-z��yY;����2�H�2 ��բ��Z�.�
��9C��|��~�����׊��� ������,���_u~����X�3���yN����ԕ5�c+ոJY��{t�}��Cɒk��	����,"�u^�{&`�ES��ڣ�I����}���x#���)�-w9���\�`�*�^������U�x,�(�B��[�w�}�8o�O��n��!�F�q x�����(Cpp1AmE�9��E��jIȾ��:Қy��c����K.����_<_��@��&P��(˲��(r�J����VԤ�(�ӈ���C	���x4�I��A��kH�CD�Id���X�C�E#�J:3&�/Z�q%��Ǘ�Rc���{��eW^����9D��k���/���l�%���&&?�0C5S��<�N^�B�����ɱ�qP'��b9u�<����9�8Q-:9p�hx,��j���gxG��+IH�m�13gy�^����]�@�/E�_�-eUE"-���|1`ݏ����4oI~�,�"Q�X{�n�߅ߣ��`��c^����sI����4?Ck����� ����Ngc��M�_� N)��=�e	0���%��!G�|S�6�(,Z����<_�a4�<aw;f���|fT�����r�G.�E�=��C1f���drvQ�UGXT "vJ�7Á�.� k�&����R����m�8��=�<���ѣ�L�����"�'k�æ�,(;�J�!�L �s΋du�]{-$�r�6��@��A�G��C,��T, f�='i�a�)`$�L�5(�R#	�"q���b��/���D��q:�GhN;&�tj�9?R�c(p)?���
,����n1��k% ��Zl��$�Ȝ��;H��.�w8�A_תI,�����ܼ_��.��k��<�ǿk����Y�k3X����k�����>��L�x�zx\���������� �����5�s���9�
�d4��|�o���ᤵ�Gh�&'`�>�(mꚣ���_�y:�&L�`>'1k��X��n˪#(��h��}2
�X���#��$�3=�_�Q�xn���11L��1�U�Ԅ�Q�gFK�H�!��fQ��QU�¨�Fc�-���4�$-B�!x��#L &�gf�2�v7�؊���:������.�IC�&�r����	;.�'�MdO����ۻ���^�߷J�,b����kò    IDATA1ӌ�TD,( d+ˠ+ҝ�n4@�!ϱ���g�%̚=O=���'J�gsK'y��X�A���;ݓ��d>;Hs��4bv>��ܠ��yl?Xݟ�Z�:������E�+pҵ�!�ϼ䑖�������siQ�㦅�MC��B �3>ȋ��z�U��[<��z)�Ō���i�����|K���;����9 ������_�;Z�*1@B��?��dA�ei�iMi���~�ZW=?րa8�ψ��+c��\</}G��~�9�YqQo�~�$LY���y�_���)�L���\�VF]�4ymd��+�?��12��f mR�#�s	�t+6�܂�'�ȧG!Z�DJQD����@8Dd�Æmj^Fޤ���<��� ��:�-(�s�%V8�v]NID&e���������gQO��gpZ�2y,d�l/�#UUg�m���5����>j�QD�,b�,g}�|�bD�A�|�-GȀɎ��A1���$�u��{к�*J1̞3�b�h��	�st��\�߹�k���$WcC�6mP81C�r��g��r��4�Z�3��bx��Km��p�	$C��\2�x�ƼV�u���d���g��|����Q�h:�3c]��bi���,&6-0��ߠ���%	F�6�y]<�����1jc�t��_�9I����6$_,_l�1�$22�Y�׿�u�s����Z/��R3�5F���/�[QQ�L�o�]�$���J\�u1����\���c�g���f˵ 4��q�2(1�:9	²��L9&�I��aj�G���ɖA�-�)Gt?�_���5����H��cH����e��0o�L��7����M0	�d�d�
�֮�3�b�.ԎD;���Ŕ�(��w��9��N��"�Cј�-���nM*���$�!baI�?A�u!�p�B>�agA���l4�d}��]��a�D�%��ېˤQW宭-�-gй<<�G���z������)U\��@W�T~���h�*�G�\�W�'�z�o ǌ��.m¾i��A�����'  �3bt�~��Ѧ�"ޛ������R���6+͛J�Gs��)�S�S����޵�h��f�w	��}�XkbYSX?#�Q&�/���;ǘ����܌8b̫��y�U�r�9
@}k��'�+
��:#���ճ��7�a��w�'��K����l��*�Z��z�x�}�!�����ƨʣ�<���K��DC��嚟�&�{Ձ��ųn�J7���g=�"3�J(9�9k�IMX )-�T^��L�@@9�r����Ap�5(��q��C���~�>''���ٺ�I�'"�DY�ǙjټC2ՓN8���,�����y�GrHF��GX�����&E�"U���G��C�A� ���g�m�H.��]{%��i)p�8�b��G1+���.����)9F�?�	j��y�1�D@����5���O�_ % �=��@Z�����{�b��"y�b�bx�C� 4|KJ��a���MJL�x�t�bX:���Jc�U:�ym�E)psSVKG(�')H�բ׳�����32�}��e��� L f��ƘL�a��/��Ȣb� �0?�Dd�g��dº����>����R!�3�j���H����Ot����";ڀ�1K=W�O@��#1�H$r�����n�#�ַq��5��ѥHj�t��sH��h-��J(�d:�db)(wPj��G@�7?5Ȋ��3M��	[��	�<f< _�^:��qmU
'��X���!(��D��>F���R�H�@8w����W�"����*����ǀ����&j0{N����6c�,���uf�UN����1����K���D��4`91�zeJ�C�����O�e-Mx��򀋭qb��3�$h�Y�(�c�͚�D��1�{qI���6�JYC�$�3�g�'SK����(V� �����3�ߡ�Y�RR�\��`l��DF�y/=R�K�b��d����\��~�z˓���x�rF�=锲$%}h}�F7?K}���63�a(�֒,��7�	��#AX�Cf}#2e�u@X���!ه��¼VE�p�@+�����z��X5�-��{�UVI�M��'vo�9�	�
s�)=���9�	�YR[��<a������;b�S�����0�]�L����vP���|M�Mz��vYǜ]�xf���֣�͵����5�Oŀ|R���E�0�m��wA��;s:��F�(
�8r�v �}dP$k���9���;��ڌ�:gfs4��"�ܽ���J(Q�F�C�z��ۏ�������q�@I��u�x�g3>�3}K7�Gm
��٬ed��0rYT���1����v0�e1b�9��tJ���'k����u7���6b���X4[� ���,�5p1hް+�*IKڈb�� t����dN�\�!��y)j@�7��	�f.V�{�Kf�Sg	�Z�҅+Mf�:5S��� ���6TW��*�z��n$6��9�Pda�Mv&���̈� O<��������W����xɊd�e"�2���j`�0&k��W]uUG%2����,��{d��X����ؖ,bޓ�
��0a~VdClT2�oai�hu�)ʗ/���z�Y�֗|�o>i�����]���~���lp�E3o�˷�	3�@XrS����v�x����Â�l3q�0���C]*@�Ў�X4�S�ZQQhkrR�̲� -�56����꾨oX�d҅ �-�-�݄L��h2���3�dA,�W۸HG_A���=)sđ�߷�*W_m)�A����j������'�����Ҏ���(����!�T}�r�T���͆�[v��MNV�z!� N�H��1c�
{~I�P1�
�z�.�b���A'3W��En<b6��8�`Դ�V���E2�� ɾ�D-�gs��|-�s��&��Z�~��YM�m,0Es��O�\9En�ǝD�����;��$�Bi���"�K a>�L��=��ö��6�(#q��Ŧ۳�Ɯ��ᕱ�}�	���4$x�R>[�6
E#�|�w�H�R�u=̲*�3j4��a��>�|�$��lvQ���0:�@�M�ϔ��b�e͊l�֌��"l�IW��V��/�7�,DD�'��}���ϜT�k�b¥0�D�A�(��A��e3EuU-�%uУ�?���H�J��H�rX4�sZQ�(��m�D�\!�=��C�G��ꋆ�� ��H�c��p!n��f��-b�bQ���؋ǋa��ߣ5)d�Z�7Q�z8����t�*M�|�Y1`�Ǥ>�|n}�,nnǀ�^hY��h�X�HU��WU,�����"[4�|��OF��� �����R\�t��i��1�`�c~�,�)�2�|�B�&�P�! H_��%'��㎎��iI ���L�U�L��uP�%8��әK��7�LXlI�?+�t��zv\�L���f]Ǟ�B��g��ڷ�$���<�A	u����l��{��A���� ��mDt�K�|#� S~��6��$KE�	�L��%]��Ra������ޞAX�`�6�bǝw����0;X�`��'�F*)�Q�����t�k���. WFW�� ���u����n-eI&�k����r���'�0�Z�ԆY������^=q�1G����@8^hÒ��5�G2Z@�o��٣c/��(��#F��xOdKI|1n�<	-�f$���������K�!�Q �Hզ��V�������=� �4�d�z��"U��d�C��G>����q�K/�1S@CMo,X� A,�h2@��|ɠ��ȡ�6)Wys����Y��-�J"��$)�D$h�*١X�LaE H�g�"��Tr��tlNx�:�E�����@�lS�"8x���#��1|���^���f>ٰ6 9}V �}�Ii�78I�E	Ѻa�[o�m�#uM%�܎��JX�F��f�=0hض(ī�s��{��A�A8D*��Ի��{o���C�TD!�6&�.R����PʛdUcq	�	l�Ŗ5f4���s����'v��|�F1V�JS��,	��P�Ed,O^&\	�����lwY��}"�췒i/���~��ğ��8wR�c���4&L.�6�:���%�ƀ~8��г�B�b+Z�A�e!⥬1������0̣�h,�S
jM�F�~��C.Z�s�b򔻱�y1��q��gMPR`̲ix�� D)(!oi��tc��>m9$��PM�:,!��S���P�GQ����x�g硵��d=7��\�R�����L{�@cƬO0�� �"$�e�E�i�I��h��?���xb�2��td�<.����c�]���`0=�%���RkQ��x겼F��S��xV�"�&`�$XW:_�=�`��tA����w�I7"t�^�9bz��kT%Sv��=�gϺ�&YK��JƐ�ŰU����2��8���=_���{�m�Y�m?3���G�rS�q�ؒ-۸C�B	�I @�!���mll�d�@(!(�dzI���EN�Ќn�V���g�������[�7�JG���^K:��=3{�-�{?�S�(�jT���$Km0j��;�i���[�����)�T�6��[��p�H��Y�Ѧ�����g�b]r���P4^i��h)��D��d��[�uB�u���2�� ��2��Xnx�b@��k�yӲFG������i�*�:�vڭ�W��s֟e�}=[�	��Qk�LYbL��U�ȲV�*�)���s��Q�������f^�<�ݣcv۷o�Fc�z��g��LN9[ъ�J#�f�Yg���bv�،��Wm�=�b�i���k[�8�Vֲ�8��Z���������3h�S-�F����6�w����A��G[Pl	�n#�G@��U�d�3'�z@C��rm9�4��A?�Ctar#t����hRć�#�ع&Z,q�8��Jb`�S ��B�)E:�9F;8������(L�}Ӗ�V��`'���g�� ?0�,0a��jZ��n3I���m�IgYr��7�1��-+l��JT5k�����'-{�v���oي<�z�9�U䈢�*�~@�RK: \���䣟d���lk6ˆ�d'���|���W�򕞶���G:0񼴷�a�ݖY7��!_Ch�u����1Wh���/��l��B�|0WB���8�p�Y��n��5�-�Yy�~kc�Y�6�Y���L��t�1*'�3Nw]V,��-'\Ӱ�����3]��ZM�R��d �d�֎�Z1!�����۱3��܊�=�vD�� Hcڦ�Bt�U��HR��+�?{�:�o����,�;8;�-b{ۭ���N���;�� D��Г,Sق(�Pk`
���h���*�H:3��}J(@b ��������
`ܔ+�a���(��)����a�Jq3���M�B�V�ݚ0���=�^��ㅯ!�o�z!=7��g���C�����$ɭ�6����R�X}��x��O:�F+��N��.�D@Q�(m[�N�l¢��nw~�VYfլe��3a䈘�R���zo�j��ѶV#��Zݝ�ĭ���XgUl�pᢧ�(����i;���B�*ڡpt�cN�7[�/6��~.�\���^���΄	Q[�}��_d���*hmIl��?�f�Ǌ��Da�y�H�(v�H�R-�E�7��DY�'����L�u3��jQ�|��#�05<|$|�����XEX��]vb��Y�=y來��l7��6�YEC�]S�Z���^9l��%vOOb�굶s|����h6�T��λ��{���#�p<@IX ��*��2ay�(̯�7��	��pi�������*��sТU�[�\�ܫ��Z(X8�)�DV2!ll�%�P����c�=�x�M�h+ŢsM�?2Lx� $wռ����m�1e�(�f޲��^Kk6�w����*ǜbc�A�`���|D����ylڶ�ل%?�7���;�*ʭ�6�ؔ�@��U�"�u��Z�8��k7���h�V�pPJ꡽�H>�l�E�Z�X��������ąLx6P�n���ƈ�,#c�s��m�4�r&�_��w&��*M�1�8H �JR-k����{�e��A���L���DE��Jkd�W ���L�[9[掙��s^l$
S�xm�E=l��;)��I#��rb��Yê��f&XےV��%�Ț�������M�׬���S^��E�Iu0�T���������1v����Ģ>�X&�H)��b�ۉj"t�AP;���0����~Z�q �$�0^U��>�~Ђq��P�ó�F�@E�1E^���LZ (|�@ AX��3�p��IN`�y�驤XSN�p(�~�?�Y~���
�iN�L�p�n���F���;��;�b@8�f�j�[W�9�@)��M;,����̏�k+Y��/�ʢ(6v�a�FMw�E�;D K��$�Z��l,����Z	�G8�e���(Е�p  <���3�X�@k܆��{A*A���|�;ߴ~���K����}��lot�����=zzk�6C�Ll��aI5�v���bbk2���H0A�x�Ҥ�t:�I���8K����7e 1��/ ��F��bma,�B�Q�g����N�%xiB�Q������#�2��ʽ����,.7 �m�V���p��y .�//�<�xFb�7���qd�8��$���#v�Lj�b����641i�ֲUa�7�'�nq���m]�Ҿ>��ݽUk�$����ε������w�i���@'��{r	��")�[��_K�l�?l��
�(YCq���tb")���&�⌹&�Z��(B_J�XA�@k��8�c��rM ��"3���9' V�c�.����yV:9��]�Ŝ��z��"���r��s: <>1j	�0��hV�]�j;��-;���[#!�0r���"����#�~�&���3ូe��I�Va������=:ك�� B�<=ȭ���hi�b�J��M�҂$�J'�g���CR\C����!g>�J��`J�	�G����u�	VI�48�8�q�g����3g$_��$�ʢ(���W_��e��󪧮ڽsc}rt�(;k��d�U��i���� �9kPiL�T��=��T:���PcQ��������I�p���|抛�(�,Ei�����\��+C�<.0-�u0�D^����ck�2S	05�`_��L,C;�K������+>i�+^]�ZϮ���ɦ������)[1=i})Y�5K���"P뵑�j[�ٿ��vgod��56�hYk
�m���A��������1��O��b�J &}�s���9C_P�A@XrD��uX'ז<!ǜ��ø���}#9���o��J�a�B
��@Mǜ����M9���&�x��yf��*�IG�� |��g��������y��Ƭ�vTV�aϾ��Gg�!�b�UXЋ�9���r��|��;�a�w�����YA�R��m�3_�԰�,C+d��� S��?~�l�+Q�#�t�<�,|���|�����2q 2.�����bb���"s�EZ a�2<��5TIN�͵��+�w��qM�cT�L� PO�37�|�O>��=Ky�y������ؽe㊬qN��0vֈ��5��&�њ���!;�<`g�X7!���r?���`N��w�k���^��luM]O�Nb;4��ϺW�����S������ߙ�Ej(N�"5����e��bLg��'~��LlX	&3�h�L-A���Ľ�!Qɬe6\1��kϜl؉��Sǧluc��r���qݲ4�
��R����=X��=�5KW���f��F�z*U��11:fqT�;����n�>icͻ԰e�#0py���{��/�jCK��`<�s��ń2�=d�jG}�~���u
�	b� �r�s�	k�Q<2 ��&��Zs�ZLx)Z�Ϊ眹��䞞>K�G4��k��7�m�ն��Z�l�>h≉� B�*x[Lzs�ik�qK������_�a�+B    IDAT:ά�Lx���.�
��y�c�ѕ�(�q���\"�]�2���L�tiG�!]Gc8�e����g��RҖ�<�'��3���G��0Bf#�r��ƪ+�xU�6,��kHW"��-�c� ��`�9�.Ϫ�'�_Z��o-+��Ʒ<}�ևoYg�4[3��*mt��ƛ�6�r�w�8��}��	D�p��aC�J(�W�dV0������En>��shl�I��ƕ'�c�NM8�����:&�âZ���2��yf5�s-�w�Ee�����8�/@�-k��������<�j�bY��n6�Iw@�՛X�J��C1j�6�vB���	[9M_��Yw�fy�I�j���j�eՐ}�?���m�g��pD��(���^�!;K#��]w�=�����!��Ć���;��X`X�'lsZ:�"#�%-�0�r����s/��:�/9��o�y��&�D�$��!˓#�+:Bm��<����WY:�p�U+�r�M�ŝ��l��$���yVԥ��=QݶWW��g�o���6�5��}�0�p��r&����6v׷mMlVO�	�V�p��I�ZRK<��,I��9B�/fZ��j8�$H,�I����T���F�2��!��31z��1NȘ�KV�|f,���
��(8¸;t,Ϣ�x��1a�; ��8�.�A���1w�7��ۧ�z��B�~>/�Wmߺq�=s6�%Ӫ)�vf���ο�v��s<�3�"N:_� �י�Hc0�y��MHb8:^�N ��_�r_� 0�I�ɤB��%��ΗY�Ux�FaPc��i� �@z��ib|��ꕒ�Y��u ` 0�zp��9���{ՙ�0/t0IRL!�D=P���P�E�q�Z�e���(�ά��6����q��N�b;zt�V����ܹ7��"u��V�j#q����G��p����nzl)1�+�\~ ����羻|��.3�A�5�e�p�$=�A�R&�,�V�VR���h�0i~�@!�HÄ�@Ӷ���9�c! sK�~�P�8TB	Yk��X�@DdA�SCLXKOq�L`b��)��n�f�Ln����B�Z�z�e͆ō�����ڨUmGm��~�y�>�D��;�x����<ށZH������6qwᘫ�g<:u)��@f#���d��#3>oD���n���]�նZ��8u��\%iHㆶ
��5O��c��}�o_��/~���\���}�+_��~����N�*���T����¤.R�T$���*�B�,�|��jn�xd���7�p��.+?��o�ڑG6V���'���i�0L��S��_~�m|t���>/����>���19�ƈ��Y��>`U�+�6(c/zы�)��G��e�]�E]�������*3J%�h4�<��I^�:#�2׿�,*?�9l�� ���֜�4K�V�&�jN�X��
Ḻϕ܁עj'�|�#�^�Ɏ�[���n�z�)�@A�Z�;J(��<@��8��Jl��{�Ln��96i�hR|���fI'�8��Zݶ��m�����F��A�k�SO_�;����B���N�Lfm��b���e *���{���߀%�(*|M�H *G�E�����9��9��7,,-Қ�_�V&�駟�u�x|�,&l��(�M ��ϸw@�	��Z���!'�8�:���d��C�Y�6rWR$k G��i�*��k5��-����xT��a[s�k��X��P��RƓWHB��2[�OYv���]�)@8���̤3�F;wn7��q*�t�Z�f��Z�W�#���!�VO[sjW����_���ojk��f����ox�k� -5G Vj���L����m޼�ﻛ ҟl��6i�3@��f�ݒ��?�	x^���Y�X�p�e��n��e�5����[��
��v�QG���?r���w��o-��{;,��W?5�UޏI�C���(���(]��X�^���yN;�E4>�b&�����B���U0�7�Zq�p�6B�2�bxp��^�[�j��֌բ�Fwo�tf�z��5S�	(N��׏�#��_�j�U{V�>s�nY\�ѱ	V�zO�)�ӍbK���8d�,��
�+�<ڵ۞2cvR�׎�lZ}|�b�����H4-gq���ց��f2������Bz{|_;j�o������% ���X��i����l8F82���Ԏ��+��\e�J_�0�BU��b.���{ca��6kr��z�#��Jh�,�b9>a���l �ǜ�qó;#$��i�B�pʚyX�ӟq��F�аM�O�Ӭ(�Z�I�؞dȎ:�\��z�M��m
*��E�G�,JS�6m�w�n{��^'� \DG����r멱04,�&V���i��}���<��x6��H��L��]N�l�7~�7|�-��E�J@ZEj�[,��_z�.�^1�A�w�ĩ�'`c��������Y0CkJV��Kƍ�+�2�@̳R���"�Jy�EѦ���=oYv^���[VX�l�S��s�s�=�%��w��_���Y���		�0��L+���xp@g
��AC2�1���a�����}��C��9��h����Š��`>��a�l�]z��G���/�'���&���q�͌�X_5���������C�En��cK�VZ�w��9�ҨϲJ�mٺ��vl��`ș�4�d� �}a@ވ�	��;fϬ���k���������ӹ��"���Jl�(��������^m;v�q�kR;��f�w//L�'֣	"�U�}'���[d�hb��É&&$`���'��	�д-�v�0�K��5fd��J�P�eq]�h!���a|1>���&���Ҹ!I�()|d^����p�96^�hj�8��{��W�cםg���)���L�2�"�-�2�[v�7��v��CF�JɄ��[����'���S�̼��I��r���g{�lUʣ�� J �:�SI��A������O(,���bA�ve�/��kQ`�,���2!�n�G�w��#����y�+�����uñ/i�-��<��[n�ſ;��Zqo��޺� �&�r�#W歳(̀���+m`u�}�;���W��a��d����Lh|4���Я�6��)��P��.�*�'�U��?�4���ц��|zp̙��:�T�V%޹�Y++6���^i�}��OY_���b���ZV#<��"��`E�,i�YT�V�g���6t�S�	�}�m�۴i�kp}�U?�A�>��ĥ�I8{ r#ʭ��cy�i�Ql�񫯲��,I3�խ�h�C��FaS��Ib?ٺ�>�7_�Q�SkuOÆ�T������r�䢋��O����ov�e�+>@S&?�$&JOz˖�v�Z5!�N�<���Pp=��U_jr�R�0��~ ���|.0��%	�����31D{hR
�%o�����H��zv�AD�_��0{�|��S�*���l�ն.��N9�,�)� �@�"k٪,��އ�����o��ﱆR�0�"�O��S�b�؉	vN<�?��Y������7�f.���~�ɳ�|��ޞ�J�ô/ɋ7ݏ@=��5��7J�^y�΀a���W� _|����Ӯ3|���4��}��?A�+-6�2��"b9���X�`��?g�@�Y�J*�[n|���� L��ac[7�&F�A�t�;�^��+m��#��;~�����(:����3(L7U�X��ѐ8�ІE�FD�{��^��0� ����]t�ׇ����+71�@b&ZqC����o�Z'�b���H���׾�56�_��9a�q�vo�w[o԰zJ�Vj-*�Q!")UL�v\���[uh��}�5}��^{x�N���M���E,1��AQ��zl�G��qbc���]��W�ꕫ��V�p_m�\�E�-����s���s_��MLO���a��ٕ!q�6��"��9���?�R�ir1�Y@5�Hb�$��N���`�i	`��@��� �P؟�����LL@���/�R��f�x���*$�iBr�7�����P�ǽh�`�`�!��E@4S�5�,��Tg�����}bi��.���l��ô�
Ql��X�S�ǿ������bl�n���.��-X|faYF\w!�M8&^�s�C��������r) �͸a�9�?2�{ �ō>`<�7�^��=��p���M>%�@�s�0�9xE8.��x�,li!4�j喛��ۖ�׌nEv&c�Y�<�^���m߻�v�O��-�='��	;
C�ԑ|���ʢ�����'?�4�������C����װ㗼�%�z�������WZ�
�I� �k_w���,jOZ_Դ�[���3�,oY���WN����.�78�i֎�����m㭛mz.kΖ �a�Ԟ-ct�I�{ѡQ��e/��׮-*��5o�^ �ÌjUkf�=�Ӈ���w�w|�������0��OHL@&b�F���߀_ ,p-ڭH�`p�4%��Ľ�ó^��	�Ra.��0����ώ]+�HzF]G��k3I s�0�j�r4�Pa�R�`�O���-a#���cR}�A�>i�ܷ&9@����������j��6�(,��Ͽ��F��`X����	5qa*;[����}�KvםŶS|�K!!x��$��\ �yC�Qʲ[�AX}�O1ae>���L�s���H�ā�ik�,������Ɲ�7c#S�`���i�a<�	��5|�w3oX�q�M�ZZ�$���׽{y�0s�[޴*J�z�}v�ΰ�/��~t������Z��0/V,4��ix
@�B+6�0 h:�������h<4�0e�yp&:�R�Ť�o
KÀ<ڠ�-��R��e��j'�NF;0�g���W��@ݬ1a}����齖M���j��r�mO)�=��Mm�aFT��/v[>�ֈ������#�3�.G(O$�lM����	�31�/8�<[�r�O�Z\+��)Mo�x5Ҷm۹�n���695U��E������	�~'�|��4O7(3��7���a��'&$읶���/Vǳq-�$\[{d�v����=�هLD�Tߊ� ��������sM�	��XV���Ua���!2�CV��@ L��D���}�z�^CB �~�m�u*���*#�������I�:ŭ
^$���ʨ�<���۾ioy���2�C�`6f�O1aL�n�%��d.�{@��B9��º�����M>!��,�ZHO�Ї܊�8=;�#9��4Db��z����g�a�ϸg�k����/
�ݺ}���fd��w����6,_��#�<�ЦU�n�iLu@��+.�0��V`1at~W�Q8x�O|��	 k�Ya	�E`R���/v�ba1���\@��]8K�9�8����u���V�,jLXo���	WҦ�F�+��<59��F��_���Ҹ�ޱ�6}�3%Sͪ��@��͂	�l���SE�U+�}�+
Lګ�� �9,j�T
5���ωC�V�l=�pk��*q��Ԏ\SN�d����3�8Ma�:`T&c��,_z):.\��59��2F�L��Ư��1�c���Ɛ@T��1S����!��$�;iC�_1M}�x�Ox_YWb��a|b��O	-D��g��j��	Ÿ2&t�.��-��νV��-C�_	w[V�H���ń�����aڌ���:Y�a�� �d\ >K�v�%k��
4��|�!t|���j/@�fQ�V|/�@���c�nYv>��p�ѣ�l���l ��pʱ'��_�2�#��.�?ǔ�I��!�#@�ae�sF�&���ԧ>�lW&.ǱZ��ot�x��������W���>A?򑏸�,P�х �s9�y��)X�<4�o�{�ڪ�ׄ{��3a4as��Äٷ���គ�c.��n����mőO��#;v��[?�ż)��p�	�Lt��� �Yy�Y�t~�@���s\j�r^4�g\s�]p�|�l9�rϚ�j��ݤ���`j�#�qM�E}*kF�mh���� �q�Z�E
�C���|��o�/���5���u���$����p����I�P��2?�ǋ���g�M]HZ�
��X�0�Xp��pұ�R"U��+3]V���@x�L�@@X}���0a����|��@D% �<#�'�g8�y�(EhgA�|<�5\�4� 9c69B�E�!�q��!�@(G�yފ���_w�ۗU����wl����+��1k�d�yͫ��[�{?�ow̱Zs�au�&��V"����F 5zaj����@f%�-˩�b���qڠ��Z�tP>+�+��a��q���Wmh��)뭴lǖ�,)@��o�ʆ�"��� 4r� �n=��Ӭ���D�u��u�glz� 5��o8��{ͤSYɒ��{�ܑ操h�>~�E���K'���U��W�(4dXb���sorӳ0����Ҁ;�rɆ�������^}�1��NOw�:�Ȕ���p�$	z-�2C��!h3f����P:�:z6@͙f�8$���P���"8� ѢP��]G���i�Lu"��!)��j�7�T���(U4bҘ���q�X��E;������4a->r��Mń���&y?�#�����4a-���M=����N�ue�9�܀#֢ȹC�~%>WʱH
 ��S�� i���p� �D��=�E�d�j�z˲���+޲y���%D��=C��W��z�k�����5�a�@�ۈF��Qd:��P��TMڏwS��u�Nۮ5��q<l�kʘ�M@ŵ�4[r��pֲ��~{��^cCu���V�R�������Z-J���A#1�%�=�Ȟ�,�)�^���a�ꈧZ�j�Zݶ���L� �g�h�ζJ��:@�v"�j[S��平&K�X�5Q	.c��}�q1MڃDwv� �C"C;�m!���dR��@N]�),g��_��~
� B�T��7�K'��hu�"#6%G��s����X��� 8�F�PH�>K��؇7��ߴ�X��D@���;�̘�Á^�<"����zO����e5�m	������3��� X�c.4�Ŧ�A����|�#ǜ@X�,
]{� ��[__gh�n�ǰ/%)��V������lN.�u����P��~�2qÅ����>��4M�7�x�[���O���C�����t 4�f�yϻ�.�������'k���e�,/nN�U7@� 4���̀&��<MT~�L���|Ql�L��W���Nȑ:[����V���?蓂���<�.��|{�S��;ئ�I�ڻ�c7L�R�<|�)\���Fq͒Z�E�~[uؓ��/{��s��w�u��~�h��v�ffx�a@T��$|��#T�M �-)����ZB�u2���\���y�P:'dܳ�е:��s��_��^/��K�!����Z����Y��X�B��sHz��bބ㑬:K�`�ra^J:�3@�^�x�����U�_h�.�M
g�B$��H�S"��o@����c �*�\��9�ƊC�6`�UeG�\IE�0E���A��_�Ӑߡ,�馛n�j�Ax�O7�Ό#GD��TQ;��g�%�t��{����;;���sS�):A+4��F6��j�@k�db<�[���T��*���H����>����B ��Ť݉�ʊ]*�w<I����nN[N	 1kY�R8S�{.�+�����Ψ��Z;K�V�əF�h�P����1E=� �uO�0���J�G.y���o���ŒP�����<��7N��~ ��|-|�\�o#��ZES.����4�	���_$:��%�%q��x���g�TVQ!��3��z��\t�ԅ�d_�H��/D551}q�N��L1S�E�EDa��3�2)e=��+W�k�cX�<#�O.T֕�E�7�����e-�^�w�����s��{�����U����֝b�^~�mߺ����d�bt;*$�����y���`�$|�< �)�H���f(z��>�1�
�g�h5J�����&���)_���l�AW~�`    IDAT�d����j������JU����b��)Oi��B�����1�Ez�I͊�d�N4ݟ����췀S����r~��&�;�ׇ��������Z~��@�쁞?_�?>+,����H����^���C e�IǗ�S@�q�����G��F-0���_j�b��f�V� �A��3��y�	��_��_v���)A�$~!�D��z�~$e*� قci^�K8���H!�'B��k���S�_�� ·�����ea��_�{��3��R� M8����	§�r����}���ǃ�)�W�It,l��A��8�b`��e����ωF���O�,2������ � (�=��P9w:�
��^Zi��%[8QO�}�<5�C�e�d�:�_�}���iR g� �׃vH�E����g��dL����u�`;b:� �{|vG�(�н�K a�L����?t��h���<�s���s��/����|����)��s5�B��W��.�[> �:�^�+�� E�=
�7rȨ%;Y��U|HDE��983'e�s����j����M%9���sN�#����i'ji!LӂT�1w�5�\�;g�yfQ�j��y�	;��~�P{fC�5ת=.GP_��5�~�Q���s�SN�`����U$��A��4
� N
'��F�q��ly�a�46���פ���~�������=��"��wz��4
����=e�I��*kC{s�����Yg��"[V[����)}0��m�`�Ԙ��n�b����� \<�����QW �>&�;&٣��r�	;_݈E��C��X�a怀Q��T�m�C�C�P�_�'s��v�ii�w��4����&���,���Y0V�b?���|���T� �H�BG� ϊ�8cpGa�r�GH�X�+"4��p���:�)�~P@x�����ҙeI���@��Ɔeնo8<��AX���(L�7�,K����1JĔ�C�`�rX����Z�ل�:�94���C������i�-d��oy�T�V��L3��)w�%X+��v �b�{^x�=�+���
zSP��3 �`,>��q�k=tt2i��7T��ھ. `>J��ޢ�K()�ό������<O����y���@X��,kS�$cO&{�a���V�I|̓Ї�9�<�$�9;[�-L����-���:\,n�Lt^x�����l->
���/JI��K ��C)�R���s�vl���t�<��O��]���eg����4М:�ZK��L����#���# �f��:�02�r��� ��G���W�)�Rv��,�.	 �zj�)�� �`�P�J@)�X��\��xY��öju׆�S�ʫP�����͢�O���J�I��;�*k(��������-��d('�&��i'C�ܩYϠ�JY:KgW�y����`0����"x0�m�k��[���~�Y�k��֣#gB�f��s�CPS"�%�N���;�$tg�q�:��clUa���w�+ic!'�AH��W_�q *�P�x�F����|� ý��k.�� ��Y`�V(�
CS vpK�=�Vj��<��������:�n�kL<7���w�(k6����^kΰ�4���*�m�i:��������H���@�@N=u�_ܯ)yL9&�]ך��\۵ȣ<`-�+O�(Aد�2��������F��)���:c`�e/!YDphq�-h\�-�/�z6քS�5��ɚ���kM�\k�I�x�n��~ޅ@b��Y~���х�ʅw��ShZ7!q?F�-T/�c���V��\Q��0T�g%��:�LXm�X�:�[ S�B1�Pn��h�\.�2,�S�V�d����"<�,�k��J��x��#��d"��)�
���kkY�������5;�nn�<9B�y1�=��|p_��lN@��Z!�٭�vj�e� u\��l:�R��_;OMݹ�N�n�u�ɱ�{�u��E�t���@��������r����5�">��н`jᙏHB	�ٚ�\��	�J9����hC��)� Kh����Gֵ�g;t�8��n�� ԭ�@�����T�� ̖��\s͛��	�����z�C���3�/Ą���k�-t�RL�C�Pj�'V�5�Ckx.��^;�����>Gy�X&\�T>{��W�� ����ڍ��U�L:��"���֥�n�^��r�C�j�C-��jEO��s���BdO�5�nv<_��:I��]{�o:�3v.����?����U��mj�\81���\�B��9���>t̡8�O�Av!@},�.�J��k���7� \*���U$���5��n��bq!yb1�8t̡8�O��Ɠ�������#� ����Aᕻ��2�:����l���2�����x\��C�j�C-���c)g.Ĥg#��ß;�r�� <��vk-!�.���5�!Mx)C�б�Z������n�Z�.�Z�Ơŀ}x�0C7I��_{�o\V9�舵;��35vA�'TMLZԂ�X3���D���d��nN�<�VP��UP�c�����	���-�U%I�|�z��}��Đ'�P\���L�ӱ9�%jf���ۻ�W�����Sx�f��y�����w�p�({��4�J;����u]�s���m�v;���<݁F/i�+����Z܇>���ؗ�Z$�����X��<%�h�������V8ǦiJ��篹�7.ktsk~pc�����6����ay�0����w	h�:;'(B�1��<��=kH���X�Ұd�i�p���� �G��8O�ε�����jd�a������S�49B���Q���I��2E��$J�����!lS��HR�}j�nֱ��:�¸P�(G�����*�	STM���+m��?�P�z�i���3�ɭ�.k��'�ND��Ͼ��|Ӳ��\�cۦ��q�AiF���3���yl5�ޥ�Q���\@W�Ȁ$����	�_����Tǆ)�4�R�<�&F����C��Ɂ0���r63.�䳁����ͬT} �0�N-c���Rjm7�	t�b��\��Z���|L����3��c�2�4�*L�Vv,��wҭ��®�WY�*��(�X5�9�td!/��|�6����иA(�!���~�0{�� <q�EY�VD���KYR����P��njS.��ԏ��7LcQ���q_�ܥ���k�K��򷵚u�
���TUb����m.���}���w��!����R��{������)�R�J8�BY��e�،,�pﱥ����X��݄�6`Nt��`57���X�Z���2a6V��v<P&���*�V���9,F��z/Q�)T$i�e�$�Q;�RQ0��ƠԢ ����UyOڳ�:[�eY�$��馛޼������9f���[�ugsa/e	�5��&\Mjv�	'y�3�+�h�Q���:p�S)e,yHm����:�i�IA �F����W\��Qb�F���O�a�}�3X~Q�	'�lZ�B�;�.!�����􋙨2�Y�a23�AX ���,Qas��i=�PLU����'��)|ń�
�<,��f-��+sB�E0lc��B�R��\����s�����t[=(�h\h�ƾ�����,p��z�v䡶�dRmH�ߜ/��a�����K.q�e)i�7�|�o-+����{��-mN"��f�3�4m{���/�~�g�����������F�K=8�9پ���x0X�W+KI��^��Wzaw�
�u��h��?��?�5!l^TB�^l��"�ʂ�	�Xf,p R45��-�P��<��� �S�Zf����*D�E�� I�~�U�:;Gk�w��$�¶�%2�(��%�} ��Rd�g�x�>v�ئ��`��!�9q�I��/��S�}˖-N� �b�c�	
�����n�+�qmI����R�禛n��e�ön�4؜��eq��5�v�e�k��ēO����η�Gn�X; ̍�TXj��P����#O�` �V&�����~�zc�e���0c���a0����9�r<�
����O�	=׽w�2Q�Ye�a��	���4������K���^ĀB=����c�'�"+�;�B@���b��H��ؖ���v�0�  aɀn���l�k(��K�K�'�`�<'8"�J�jW9� i��9��]��0hD[i�����Gb� �oj�K,�v	¿�� |�o^���M���Rl�C�ZGv�i��/�ܲvn<��x���29U�Rab�00d�*�.+<��/~�M/��<�����њ�~ɁƋ�n�wgl7�=��-e��e-N�(*�jgb��ahW/�ζ�8���Ga䅊sk[�wo�7��"�p_1���bcQ�����W���Q�Z�F�� ����9�m�v3"iv2��eIKܩX?_�I��g�1t�! L��"�0��7�W��fN!��ga�Ȭ ����Q�I[�I��֡���6\��5{�o���k1��"a�C;�l`�!��De�7��,���� �]t�c��,���.�j�	8H��l��?��[c��ҡ�<o�q|��7�������9/� y>��ڵ��K_�[�z����?��[������&+�#�ѓ���D������V/�3Iit��Fg�O9���/������c����ڹ�^���l7,Kؠ(�8�,ɫS'9N,�k�N�V��_�E��/F��,�V��hP��;)�^l���Y��>�������J�e��[�1ױѴ�Z���zll�iQ��r�FjOY���le688�+8���B�Q&S���;��X� �U̖��3������|��*}�]R�F��u�O9>�n��\�(��Śb5�0��{-{��?V��BKAE�`xX~�0m.F�lS�������}!?	�ɑ��o 5��O�=�k�����~�U<����E�����pa]*s.;���u�s��8������}C����|�+�|����d�&�gc4 T_�9�[q��
sN>�dg����q=��q��c��o�j�A��m��	;W��k��֝e�{��ܽ���~���*6�,�]���[f+���I�1!Y��h�dx(�>�����4 �\���x�w��M��{��^�A 4�Y8:"��͞�YO�~B�z6�h�������f��a��Z�����e6lY�kI\3��i�a�5��a�Yb�%Va�O���l�;.ge�b����Gj'��am�f�eyϰ�6sKz��m��3V�V��L-����me�ϵ�a�X��ڛ�u���y��Ō$7	D���x�ٖ��arL46�\�������w�f��ª�������Ҕ!&��K.�ĉ�fѣ?'�����I���/�r�s.s�c�$,��ER���/Ӿ[c^�G[0v���7� �@���`�� ��	�8�GO�,#k�~9W�5I"�"��M�[`�ӱC�g?�Y�GinEQԊ�x�7���SO=ud����6��8��<�ЦYk{��f`�����?m��v�~Ӧ'g|�L^�'l�':�	��ɁHs�I'������}��a�	X���Vt�� bP�����X��Ă�[y�jQ��<��x��8q�L:I(l�Z֞�a��ڶ�/����G�bGyӲxڢ�U���ȗ��;9�EHiɄ�J�;�K�]�YT+wp�,NSk�UK����F4dI��%�j��Q{�I��'��| �PA�.E�ȡ!�L:$MS�R%�cذa�O\,��ǒ�<�����k��a�/"�"�gԜa�/�C&.��s�)M�A��4a���:�|ļ��gø�a��Q����a�.spbΪ��	�L 9N}"�N?�tw�}���������5�\�D?c�FB��� �Cb�8�5H m#�!��̡{�<�c�����]�& |�5׼���~��e�y�sS�3����f�x��m�5f߸�߭VA̮�ꊼ�nv�VEn�P2�:O��@`�������?��yq ��
�x=�Cg3�B��x���0{�r׮7�*���XiIT)w��,�&�'��<֞s�����tݢ�bI��X\mZ�'���w�d�	}cP�� �Q,X9{����\��l��&����V����rа�9�k�������oج�Y� Xd,�tJ@�6�G�,Ą������A{k��<y�e"��_�җ<tJ`�6 �r�).p�o~��@g�}�?; Ä5��k@�� uM�����jC9 ��cN��\r�ƽ��Z �|G�N��W��Ua2��|��׿��w�
�q��	'�`�_~yg�^���9���'�"�n���e�6����9����	(�T;��L𓍇_��W��iG�{L��5��`�sЀ5Ƙ[�c�e��������V�Z�Ե�^�{�
�a�p�^q>�����Ͽ��z��y��=c��o��v\�E�C�����n'��X��:�,w�}�_p@�e aJ��c�a�p [@����$Q�\�.�b�f��Ȧ�Ik�T���m��
���X%���l������c�lz�NK'
�7A��,�iY�`Ū�Ŷ���<~�[�ю����۶�ڝc҈ݛ娋͢�5�A�6�o���-�eo͒��f�8lV3��C���x~&m*�!dG�i���g�s�1�MXk)�MLv �2�9�Iʀ���w0Pq��9��#�}^���o�������	�L�߹��s~@X���Ó�1��&���#X��� E�m�{X�|�V�d9���-&�pB���SR	�ym�� 2t LX�ĵ�8�3�]v�[ь�?��?��(9N>(�	��/~�k��E�v΃ �lն�Ap��6�m�G`Hj��ԧlb���J��'�s��o_V9^�{Ǧ���s�� c���^l�}�y����۶<�S�Z���+��C�0aq ����!�����eT�kݺu��7���$�$���4 �Xߩ pX��l²Jd�z�=�����ZOo��m�Ѵ�c�p�����Ǝ�Vi�]�h5'-%���e}+�ĖEm�-�=��� ��P�x� a�$��u�2��5sL�Ul:^a3=O����f��Y;^m֬����Ծ�w_qYFN-|b�1a&&�����ĵCY)���B��cp"-�ޘ��������W��c]ˮ�5���������7��#cx� ,тL���1��$'�m��r�s�m�	�9b�!�s>}���w+����˄�L��/���}z��9c��b���+�饗:s_�YI�	$M���h���cq��8H#��c�>>�<o�qr����o۰aÞ�X[���>y��G64��E&*��u���_d���o�O~��U��E�1�r��蚼2_���,ei|��4�-���%F������J�ַ��l���R#�CL�*+W|��
p-�Y�ֶ,�,�*����v�ŗ���g-��m0�a���,�u�ٞ]MU,��Fl�hOZ�3c����-�"l� ��ٝ� a�+�S�*�-ɩ��g�����E=6��ht����Y���hX-��*�c�6����_g���X�&�b�0Z;�-�`��F�H�?�2���!ib��hh�qMm)�?�'V�&�R���X��Zlh'_����Br����Tp b.(K�$�D�Lr_h)Ѿ�'��C�"�\���C��9�(��a��ǜ��"�@�`�,��]���Iý �<�^��Q�;�ڗş�Xg�{���CF�P��p�m߹C�ҵ�(���k������]Kc��ʇ�l^i�s	�":��O����W�w���>K[ W⃆���$E�<�< Ecȁ�g���̅�i0���I�~�s��f��s_:�L	9����5
 ��v �����s
�)���9b��N�O�g���X2�ǲ1<f�j�5�զ�oUb����q�2L��H���V8�J�!�'{��t�&z�x�{l��j���#,<����md���zWZ�ƶm�öi�-�Js��2���N�ðhO��2@��(�+�n��̄�[̈́T�<��O}JP��d���?}�R@�c�J�pѓ����R�,�қ5OȒ��EVćc`��0����&/?O� }�3oC�l    IDAT|�j�p��a���_��_qf/�<c0&�a�������>5�Y�9+�Ϲ9�p>bi�=��},�x�y�Ґ,­۷�5�$i%�ʧ����߾�䓗�	�����գ[nퟙ<��nX_������Wٖ����A��乯PԐ�a���D&l�N�� ^:�ق�K���t:�@��y0)^���q���| �55�+�eI�</��9�γ�/�Ģ���̢�n��X��n����{���VV��U��5,�N��a5��Z֎�;��!I�j�p�� �e���{F�<�i"��L���DGZ:t�eC�ۤYd5��j;vm��}�c>xh7M"9xfs̩M�,&#�KE1����4�n��IqL(h҇�-�&� +[I�|6'�OZ�9�&r��������=�dԢ���#�����R����ʜV"�/�*�G��:�#s&�~+*�>Ww{� �w�Gڡ|:��=��7֏�p�6�关��q� �w������cz3DNl��E/z�;���	<P;s/$v�`c��"cY�q�ߐF�S�Y>g����_�ӟ��M�L�m�I�r����v�o����G��:�Μ�8�U}+�5�y��+���g�j4Z�P�xb�$�j���x0Y���á�`��������x�
N�����c�G3ؔ%#`�SsLK3��YVi9�ҺmX��.��R�)�Jjq{��{,�����Z6�����*�%V�v:cV���ê�ͨQ������ a_�<��@���C����fU��W�Ht����[{�6c��y�؎];PX,�����^����!:�1x?X �-������\d!���A,	-��_AցE�,��O A��<���m�8�o �v��x���с������~�/H z@�����':��G���x���G?��Ge�2��_���:I@� 7�����d	@�R�3�����I!�$�3Y��8N6�|�o]�d@xŎ��4��#�VWM{���8�t��o����5� ,�S���LQ�w��*i�����/ o�V8��I"a �)���/t3X�k� 7��!��{��k�P���t'-���ε�/��(Z�T2��^�w[4z��'�u&� �V���X;�*@xM͢����aq5�v	��Q�`����펼*���DByP�ØV���Z��K�i����Q�,J|�	�s�T�ik@�I:��B5���̈́+z�@�����2�q�2a`8|��$�[lsR����
��b�k�qA*��s ��b�1�áDԊ<�rl��cɄCfͽu3aƗ�Z�Ҧ��7��1�7n��G;]u�U��}���Xrh ���'���'|&'��QV���NEf���yqέ��Z�ǝ]N�8�6���w^��������j��;o�=�R�#�Fn�x����r��{k��ۿc{��u�T��<�FiHҠ��cN|�;���d^�9A#6��/��l����'��AJ�22�^ �=�q��(`^;����n�;�.-A8F1Ha»-�{��L�rĄYҮX-��c�%�yâZD?��@�9Ⱥ�� �Y+�!�c.+�
��ؒw�5�NV�H�p6�D�]{v;v��qhƲ�	�	��e�jA{����-
c��o��+�`EL�4j�έ��q  YʄY걡�p+�S�E���X�򗐀�sa��_���X�ɯ盭m�N?/9B�7�q� �u�n��O���6,�$0��?�tX+�p�X����q��״��44?���tb�C_@���/��R�7iǟ���w��noodsc�<@���e�{7<�l���n����L1xJ�`Ő�%�=7Xw�q^ד�)�ê"ݏ��Ӈ?�Y�t�M�'�h�l�'g _��>�B�T�%B��l(����S�f�����B��jn��a�#��,۽���أ#`�E%Nz� Ѱ
L8M]�)4�"Y�x�Cj0����d�I9��������׃ӡg�4 l5��9��>�яt������t>��оfa�c�	˯�s�Q��I$����d�md<���BR	��c	�|� J���XwH�[�O?��uc*S����Eb���ǚ	�ϸ�L������w�	kH�j�P��i+B\�z/�g�+	��"��t/�"p�9VQ"�M�0�JQRT9�r��]{���}��q��y���Q���P�jN3���U���/�c��ۻw�'+��t`~j��0����d��<���48C� F������Tx	�F�����A<���`Z��c��#�~~5�ن��y(�9@8j�#��{��=�-3���,A����6c+V�XқZ�Z�	�{Z2�C�ps����,f�T�פ��4�Y#^i{��>��Ԧ��1%�k�}���T�͹Js1a@9��	?� ̽�AĠ'.���������cG�C��c`���`�9�T��}|��G�3�I8�]8� a�5!�<�����_�LD%�������!��� bƳkLз|/Y� #sN�j�n k�L�B!���q"|�aI�\�q���u�D��Dj���y�F�����~k�Ax՞�n�Z�o�Y�*_�o�y��G�e�\nO}��;&<������(�a�_q�����XB�-��D�������;5�u�D�|�΄��S��>�U�2�(����b� �ǹE0�ֈ�,Ax`�f��[2n�kWc���ZeƆ��&��N����v�.�o=羞�QTS#"���URSw	WJM�hOk�LM��Շ>��t�9��҄CGR8�5��ßgt����,�)�i�L�C,1$
�0�1@VĠ���9� 	�Ysį��x.2�p��_p����/�Y]�7>X�9�[��$k��m�I{i�S,�p�=�UD6�X�)�X�)�_�D�(� ���H��e�b���gL%I�믿�ͧ�vZ�f��W.B���?3���6��!k����#���ϿЫ�T�&	Ńk�X�y`�[<�8�4�@�QQvV:�A�7�/`��8��C�r����}��sˑ����9b�q�!e0W�#.��b7�Jdyk�V$;�2r��>`�.�plQV�V%����:m+�L�A&L�Kg�D�)mY@[�����F%6�䊈	��	Q��m$:ڲAs'�t6XD]X�Μ}�`�s9$�c�b����v�-Ą�cN��B��h�D_�rR�����B�L=͇n=u!Ki��h���}bZ�З��u2��C�gZ$�Gat�Ƶȅ���d�z���&|�SV��WI�q��9a���r��>�`҄2L� Ua�*����5�/�o��^K�\ߛ$��������SNپ�q� ÄZS�Z�EloT�F���N��Xjδl��՝���Nx34�J#�aa-���.�ք'U�X��Z�X͘��A�j*�.!}�L8�T-w/<�#S�p�:���+<�"�T��{lE���?���,ߵ�*�5/{�&�5r�iZ�cվ��6eq�>w��Җ�+�sA��je��q\��OY��cʆlĞb6|���������d������G?�1DZ�d��jr�=4i�R���sK�q:<<f���Xf�&�)m��	� e*�1�m�p�R3��g�1ǘ����l8)�pqYʄY�cgc�ZS��-+�]�q��r̅���sR>�;��?m���e�"�[9k�gQ�V���\EbѶS�1�P{�f��o�qE��0[,&$Q�^�B �(�`�~`A��$�Y��9�ƊA��P�?n�⁤�J4g���r6h@i i ���x脜�/%L$��#�4�(���iIԴ���%�\ayT�(�ytĊ������F�|�KƫV�H�Ȭ�p�C�*}��(�S�"G[^��K[�E�(k\�#��&Q$8Sʒz*�3���3,>�Z}'8[Y�~ddrY@�I���c�Q�θO0 ���zʹ�@�u�j�Q	a�j�j�9M�p⨏%K�\_s,�� ����{����\�x�ɿ\�/'��_��x
�R���n܇�Q���e���A���b�b�ݖ ��/�
#���f9ڰ���-�p��И�Y��H��2�3����2���~�-��/��/����u�-���	�\c�2�wZI�h�������Ԑ���JիÀT!l��,J�Q�7��}V�����l�����c@���V&�,��c�}�l�N�Ɖ����0��,A�m�h�ab�Ҕyw��>\�1��uΫ�!�"��|���3,[>ѦmЬҶ<�ld�1a&��61dEcU�"\h{+����<�ؔ���K�FAh:s]9ESE�/���1�!�-3�X�/��J�S,5��D���̧��a�@�9����zDu&�8�� _��cT֡p!|v���/��4~��y�RP}�ꫯ~���)���d����<�4�pjUY�����%J�����>���2�H9v� lYW-&D-�a�L���"D-�A��ȧ-�4l�0�p� Wr��,�Ȏ+�E˨A�����Sт���F�ϩ���^{�e+N�f߉6� �~��ޑ�b¬����M�y'����j cn�?Ŵ���9� �|���2���=F�_�R�Z��.�*G�sD ��e��|�X��
L����+��\[	�}��jĜ�[���	/�8�!�MC��M��h,�3�|�mY�a�yI��tssi�����v����F�đ�NTCΦ	k%�3��.�@���>$I�˄�j�~h"9� �K/�ܓ!�J��ֈ��wX4r������[gUK) ��XTi� L�ܴ���R@�eׅzV�q&iCr��QA�cW\`�$ =Ͳ�S����0���yj���oM&�IF�$t2���>X�ژ��!kcV�_&��JJç_ m�C%� F�T(1i��g��Q�D���	/��1�YHHr^��#Nrڗ>�?#�x����A����1"���>d���"�K�-/dg;&���tȴ�H�� �CK�G�<z-(:����&_z�;����g���W"��	��6�&�Tc���� �!�sp���39��%GT]�hg0��ˊ�JdI9b�%#�Z������'2KҚeq�Y�� �#T�_���˗6��w6�$�W�k�gЩ��d���FO�lų��m� �,�ѽ{��f���^�2�F�T{j�G���)9�|E�p����`�&6!�h� �����7�^�0a?���>Iԑ�|���x�\�+���0a�@E�f tZ�	i�(���8"p��
�|���x��F��6n�ܦϥ�ӧH�:Sd��R���$-��]J_���l�fr�"fb�]-�"�)ZV[qLX$ܢMU0���f�{m�j?�Q��kU	�y��р�*�P�;�,11�Q���B :"�+%gv��뼞0�I%�>+���z��l�6�ɖUҊ��m�M�jᘫ�1iqMv[TM+��[��Ow�#.�Kf�;YSLq�&�a�c,_y������h��fY��Q@���̈́e�2Y����U���r�i��M�|���5�b�3i�Ì�WIH Oz��)r  `X8p�!�(*JYv;�y��(�N��@����!X`�B`����I�� QO�0���F3>�Ѩ���o�)���`GG,��"',V�~�n��cDFĞ�\Z��`�>�/_}�տ�sg��u5��թ[��i���!u�:�������D���`��SO��CmR�G�����.����]���c[,ݽ�l��!jq^5j-��=V#m9���kl Zh�*a��j�o���L�D̡^���m��\0e���h�'Z��X���Q�3��>����4X%�҃Bט�r|Jv�x&.Z;(8^+�ˎXv�Ez�yU��3R���1�n���:Ąa�%bQdn E��`� ���N�d�J^�| Y���IW�{J�R�������S���g���.�Wu;5�ĈC|���*`�v�q^����C��F�`�c���}q�u�V��&�LZ�S����aM g�e�p]S��YAè�j���|v ���m|z�*=��f�%qfg�;�֟��B���6PkXOk���wZ��Vk�|��vj=l5?M��*=��V�ޟ[�PԽ�l7.����
�}#ϝ+I�>���~��UkE+m�~���Zk՟b�jeв��G?���zM��[�_��~�U\���M:Ҡ�6���H�..���Ċò��$�����������c.�ﰟ�]
�׸�<~��)r!F�x�<dRr|jQ�I;�a����J7�}��-����B������=Q1�$%-���{~�%�cMDI�����g�kt��>�YdOq3ܛ�l�w�Eڂ�BB�=��Ӓ��x�oX�d���4Ԟq���nMb���g�S@��0Uוϙ�ܸ�e���A\#��al����X�a����^22'.��g�L����f$��@�������ZW�hU��b��"�!�	�[���ZwHXk�U�j���T��ֺ#n,!�(��v��������͏;s���0A�>�<�ν����y��|��}�{�ѓ�jé6<���+͟�gޞW���J�f�ғ?2�������4t�})�R����fͭ��Y�)U�2���Ŏ��O��;͍.a.�p��G�s�A�[ޏTSo�i`d��뻺ӷ~�5���z�>4+oo�?0��fW�wݞ��pΧn�b�A����ٌ�Dd��@ϧ�R����ar �5�/R>s@ǙT�d��B:K�C����&N��O�y�:���s1�`��1�J�@X������0�H��m� `��;֔���˾k�5LG]���0<�L<rue�jo
ޭ�8+�3 �A9�� |�����-����h���8k�O�B5�.� ��wDo
���W�s�_5�5���R�|�Bc5>!����T��I��q@`7�����Cs����ݝ���Ҳ�H�<|ߔ�ߛ��G<YB�!
����9]����b1Fa T�h��l�+q��k:X�\�J��4R�3m������Mw����4�wn���<��I�Q�� ����YC9n2�e����HhG���mTpqq�!m�̲��g2cLؕN���;qO����xV�F�q5�u,�8(f[��j��X����`A�v�(Q�6����x�5�hg�qħRg���{%�8��?JأP�K��w�H'���1w����Q&��'�y3�ޡ	+�\\P�a�N/bt�9�����gܪ�q����1A8�Sȫt��z-k��*}i�V�	�{�7�=u�t�K�z��<�r��Й�׺rv}v���~�#�d�����0[�0.rDd�ݨî��H��oY�(r���M��J��3+�5��`eϼ�ܬ��42ܕzq*��	��;��ul;D`G������y���'׍S:�����ц�e9��x�x?l�)5�F�|����e;D�}�m�q��� %��I�siyd��c�D;����+��}G ��y����Ĉ�v�s��&��vm��x���0ʛ�m0JL>�q���:����3����4ox�ɀ0�0;k�	Ä��p�O;�y���J��p1���r�Ƒ�ϲ G%��wݑۥ�+˶L� ~��s�B��,Fm���C�eO�>�����Z���	*Sw_ޝch�Z=/ި�i��)'ú&\�z�����	�yϏTEbIi`h0�V� y,�����ޑ�T�w��=�RmhG�&�N=�p��:C��� ,��ь�6|Ɏ�%�C���dJ���#(	XN!a�q#˩v��:_)I���"HH$�t:j�x#��b�`Tn�g@��8˱�c[ęQ��9�_���t�o�{�A][�;,'��4ͥr���qF�����ׯ?���,:�m݂&��2תEn�rr ��I��ȍ��J�NI�C�C��	�����F�GϽz�w�0�#�E��0�X�Z-��HwW��3�D���ONVv�����W��9�C��v�V�'��x+���H�N��ùJ��m    IDAT�r�E<p��Q�w�``뮧
@?RO}LS=�{G�}��4������ԗ�#�4<8��K}�l4�8��٥��LB���k�Q�ߨ;�3؟�E��i���kp�ZN�}6ʍ�ow��S5`m[���R81,�6�2M���(�U������	�n�1��o,�1�Y�`�-r�a�ܡ�R�Xvن<�P4%1��` g{5�0�I��� �c �V�����	FA���W�[����a��{��-7]6���ı@�o�G�$��RHC������O������
�����n�ǘ{�D�q�T5=�c�
��@h �f�uో\�Y�������Z����,��\�I�������`���2-'>���`��]����袌"�ew���ݬLN�Yը���]i�p�W�){�9���T�	�y9��3E�����4_s��؉4���O4����S:�:8���I|ﾲAX��Fg4�Eu�������v1����m�]��x Xx%)�7�x�V�C���f�Q��Ⱥc�&[�c1me�Y6:g�D��O����a N�û��㽭�Z�FR�O�]����not�)o|̂[}ټၣ��#�,MG�<O{`�,�t)0@L�#��,����H����F� ك�կ~uf�9²��_�%}����F�lC��:t\l0�����@�DO7aa���RO_5m��K�>��ޮB��W
�2�YlW^��f��sNI9�0����bۣ"�;�,3Lf�gw�kp�t���*��ix`8�)���]��h��3Ə�k QFh�c�'W�;DD�O��9U�N�DԣǺo�X˯3���d��8/- ���h)A"z�%b���l���9^�ԁz,`�H}4c�9?ړ��l��J�2�";��C`x�@\߈+���X2L���$�'F]���稍�GA�̎���3�}�­7_6����f���������@魥�G��z���ܹ{��}�ĎJ�!���cB� 8a���I@dtTSw�[������8 ����,6d�Ҙ��[��e 娅��JA���ʷ��b��w(ݦ ���FW�!d�P���G&��.'|gq�+��n�1�sfj`���8#V��oH��t�Ȍ�-��/�F8P�q�gnԈ� �0Y��y����q222R�V�W�^����������qo��eF�����>�ꛛ����%��}.�g�����<3Z ��;zEu鄃�`h2 7	?H�c�Q�6��F$������Pl�Ɉ��h��2��t|���f6S������j@)�߉�!18@�~&���0�S��3���v�Q��0��7�*gI�3GI$��N�Wv�t�pT��U��O�Y��� |���{���n�t�T[>8ԟ*�=iN����כ�?���'<6���?L7�pS~xG&
�X�W��2��T�ёyg��I�u��(lEr�gf����hv��yի^�+��@�0vT<��L�����=k �����/��>�����ӟ�tƒ�N;-�ڏ}�c�8i��'P�p�	YZ��%��o����p���*P�o�t_&<��U*��֬Y���2a@x��o�t��m˙2�T����ZZ�|Yz����n�rC����#�2Y�:#�9�@N [�8!��lO�6��xE��9�5�C�1B>�y��K:/���V��{�}��5S�����V5 ��߮]�6˖��H(Dn����gdݖ���o�L\b��g>��!���Ȑ�W�z��椁�q-�y3 PwvF�X�j���޹��9��d�	���+_yR���M_��������<t�=��fu9�0�0
�;R@�'��e:�ta� ����f$#/8�{���8H��V=��L����Y�k�o�ƍ9���?������s�T�d��ߌp@�$�j�9���~��8j���c�0��Db!��?��$����3�Wz���z}���s�ʋ.:�裏�c"�9��Fh���vå��+�g����:��?O��vk���'��0� -q�)����lt_""m[��]ՠ��b�w[#7�|]2��f�੠�,6.��d��D*v�ؙ����� }��~�Yge�ǌ�+_�J��t�Iy{�ؗ�����~p�햸; �n�`~#���J S@��	�u$�Fd�w�'�
}�=ц��ow1�p��犕o��G�a^t+ <�"�k�w�#Z�^�����~�����s�c3� � �a6�y�o��%nh��~�s�˕�s���>7ꄓ2�u�ע!�hB��͵�1�i�0s������	�N=���p�%�4��������H� "���,�e��A3k�M+k"}�S�p�br� �W\qE�>�ឞ��^|�9aC�fo�gEo_5uwU�҃O/|����?��t�/�z�}�
�ٳ�l�~�2@�QG����k�"F/�7�q%
�d���'���m�љy��)���vr/�s��㙹�L����k��f��0�8q�� ��_�H ]�3��
p� +�~�QGe�fd�=@��dʞK@ 8�}�o����+�+֯[wnGW̱Xc��o�l������R�қ���)�9�yv���+;���B~ (M�e��Z����<������+���Y��-�tR��Db�Y0�py'ͭ����L�&w��؀+4[�4�+O�r �剋����&w���fj`�5�bR'���$�����~&h��)�a�G� 4Y��~����Z��֍�pI7�s�x��g~��[2^�j���+6���Yf��n�l~}��=��'�bɲt�q�������0�,a m�/�1!F�&L��f5���e�\�E�`ʡW�� Yco���Lu�Nfq��IE�+��d���yqE���������@���g����]Q�#��������P15Z�hq��C� +�lGb{��h����a���+s_��/��8�8�.�i�;�w�i��V*�׬^s^g�#N;瀇ܺu��{�Ȋ���i�cN'��������?�M{Ι�����a��v|+���n�v������O~2��6c�,��F$e�mres'�s��
�h���I���,Nڽ�T����u�KY16�nq��<�{Ϝ;SS���J,0��MDF�Y��=&�r��/� 4�4\���0�p�o�;���D]�w�e��&������^A�V�t_�f՚s:
¤�|ح[7Ww�Є�ki���N:���Gw��7�=�Tzs�'t���&Y�s#���k|!�Þ��?�3�ۿ�[�B ��s��:(k8� F�1`׀.e� e�;�	�G��Bx>���j��:�����['N��aДGО�#vU��\�� ��^t�EY����?�#�d����?���o0�Q b��׾6�� ��nr�{��9���H$Տ�vf��)��ȘE��QЮuww]�~��7tT&����o��{��O�ф�Y��c��yp����t�w���"��K��� OY+� A��d��J�2�&¡�4�!`�nXhs�4䪫�ʂ��J���54f hW��PN��N��v���� >S�������������vjv�]Y0^�[VŲ�����l�1c�g�}v�	�����Fg�`;��&�� ��A	��s b���I�93(�b�.�Q��bnÆgw4�;�Ϳ��s��S�v�sC���_�����$n^�|���
Q(u�Ȯ���p<������ׄ�?�ъQ��/̕�bt^� �ד��f�\	CÙpyW3�VH���it��1���u&�{̲�5�z�_��;`\^54�	O��g��d�G 
o�۳�K�6������R�>��<�Ɩe�XDz��$n �a����q�]�'�;,��C̈́�%��G��q���wt{�%����o�_�JN-�F�J�?���)G�'�����~�n�qK�XP��S��0.� ��̱_#�3� \��9DE�(X�3�1�?'��	9do�����a��"G��-o,�I�mv���D��`���@t�KYC��e���L�`�Vlذ!K���Ӻ�;F��ۿ���س)���! ( 6�G��G紤���lj�#G
������>s����y��כ�=�,jh��g�K۶ݗ�~��t�I/O{�~��~��F!e�N	F�_�# ��K:K����_�r��-�y�a�/x�r���5k�Ne��LN<��� �o�FFD0�.ӦL�>��g���ەe�i�d�Tˍ ����͙����Uf��n(��L]���`R&'��7~��,`��'V�� 1��b�[臨�p.�{ Q��#����(�����ի�\�b��v����]�����7e9��-��3��N��f��K�����G�I}�~���0��.tH�V�e)!���qn�"�������z0Ss
��%q�X 6���#x�r:$y~�ɑ�ӌ�q0������kT��1F�-����5���
����=^Wϲﭞo"���xl9,��R��~��(�Y�гo䑳��F���{�R �v1f<ΞʳJ�#H��m�M"��%쬁4qd�da��^�)���8��� *)FGv�Z�z�ʕ� ��nټ��}�u�����#��?-YrDη�*5m5��Ί
�~K�(}�m7�V��^���F�wݷ��T������Z���t�TA�rǎZ�.Q'�Af���!vJG�<��&�',؄�+!ŭ���k��xJ����ࢮ6è[[����8��Ȩ_��ٞv����a�!�dL��nx�mI��6NV�QB�OJ�F�����$���	[X� ��.���?���!��f�h�h��F��.ᅷlټ���c���]��7¦��4��������ex yHqTعy�^m�(�Ȥb��=���P1�Л�q�2Io�6IT6��ow0���pd�J�*x���A�E0��z.l��L�S��1F��-��'	S:;*���L$�re3Ze�����|Yg?��>��ːe_q`��9 ��Vl�����,��
�'���q�v�ߝ��g��]�������h6�C��|����E��o��	Q[x�-���C*���Hv�U*�y{��jW�>��R��E?!�������Kv+iTP��9��ў�q�^+�����Kc廨�L��L�}��F�)�O��m_|n;��c,c�0{����k�S+CZ�aꋲ.�tNɇ6a��3Jmۖ���3r��V'����2U�Ҏ_f��]<�w#����A�ߔ�l/�]�����S��о֭����)H&�G��ܡ3�BWRg{Q�Q��l>�jժ3:�	��޼i�4�CԈ���P��+�y�{k�l���
��x��70�w
^��G�|���]��q^�{E��4��=;�Qv�^\�5c�.q�ȭC�7"�����ĥ�tv��#�N�G:A�rQkC�f���#{��Ap:۾�{��r�38I����?���U�5/�}N-Y�ٶ�ɸ��rRԊ��(��ygJ�_�g��c�?S�֫�R��D2��,�D$���J��yΎ��[6�ڞ�p��I�ၴ=��k��OIc�Ԝ�8*;hQ�N�Ai�\S/��0��זEG`�#�*ǎ�N�@�B.�� �p3:��Og�dY�I&�(�jL��п�y������~G��҉��`��N�M�{J:t�Z��$5��Q7XW��������՚�f5�2�*)	��a����˱�M��Hg�;�	��y�������@x��n!w�15�UO��	���L8�q����O�n��4����5Em3o��:�h���ָ��8�
�ց�6�8pJ���{ �a��>��G��� ��.f�����	�'L ��� z���Q����v�{�ʜ�҇�oY�ˀ mI�	��� Sf�T�s��>��������Y�ǎ\�GR�wfBq�Jh)�%�ҁywg0�팜:�e�\g�b�����,������R���U�N�a�ڞ�ێ��Ɏ9�-��	�h��6,&��,I#��� !�Ƒ:N)��N:�1�?Fi����S��`t*HG"� ̋�ynS|�8�!lQ9��Y6��g=+k��I%�&uFAX=��pʱ��N$�)��κ0�[��e�W2 J���?=�����G�đJh&Z%[��,D`�5�g�����Z��c���S��T��0��ݩ#R�������X��uhc���|NyIሳJIbw�g�$1���sٯ��R������Z�~n�ʕ���7�ߐ#p�EM�|�lo4�+�k��>t�si�udgN�v�!��=Ǻ� [�3Q$n���;K��q�-��]�/����A\ո(&L�PLØ�u �h�>#I���eS�9"o�z�U�]7��8c�{�'rvz���������%3b��SN������75�K�_���e��o~s[^d#�"	�7� 6��~X��C�^p���X*�c�2��h��I'�@rg��g<�`Vf���vlD"!��>�6���[��OG��U0�@�ddƞ�3�,����V�^=} �(:�*v�8-K�h�3���\�� 0�����j����@
`	[24�����v��rm3�3	�x)FX��&d��> �&�S�k�0a�2jSiߩ���p~��|֡e��$a�h��?;ǰ��$A9L�A�#�Hc� [����`�.�k�\���xΣ=a��S�^�}h{ڗ�|�0�^�r�=ǐ��킢��l�ϱQ,��V}��~����ҁA����l6bV�Si�f��e����իW�:mL��
��-m���:[�L8���P��u���a�9�IX���z0 ������d(LU�6�9:*�ҹC;q䍨r�B�AnP^���7\[�w=�s�<e��� S��v����ߣגf�J��A� I�=�i���h����m~Е9����r-]~�3�%�����n�àMx"�Jy�=8�<����L���9���� 2�2�;x5g�o����,"�h�e�Fn�Kwww�A8�	�~��yC�O6:b,9����� qA�U#8����\!��P�*6B+&���Q^�̹���	�+�|yǠ	�1 c��YB�Ш�{����q a�q�kP�g̯@�W]	�DD����Sov���:�6�kE���I=�qw���EG��Xe���}۔��3 /�~�����3�5ϋ���V��
�9β웂0ύ�20�~?Q�PD[�n� �#����s<�Y�/�p3v@��rI�m�i���O���'�v�~q����oy ���*�,NכU\������@/w�����l��tZ-/?�n���~�ba6����Ɂ�@�5�N���AE9�c����܁t��=\�)@������O[I��TR��xw� �m���$�h�q���b���؆�q���oAK-U�Zߋ�t�ǁA��;�C��bߚ.K��-Gr6D��3;�)Y��r��>��������_|�i΢v����qæy��O���}F�q��fc5c�>���]��@��)_�ȷ*�n��ǁ��bGta�L��b4�XSFt?e@�Fa���D��q�n>˰"s��щ��g;gy���;�d������:���d�N�e�����`���]�F=��D�1��vv�qê<��8+⻸�7��LT0���#���a����P�Ѫ��V<>2kYh�-b��e��s�7�'~�Z�Hi�	��&|�ƍO�hRw6�\��f����@��M.�"D��м�HV���)T��+O#�M��݊I�j��{3@m��~�!�r5�������}���L�-�h�YM����0��b�ttbK��[Z�N�k��5T�G�=ֽ�S
�D@�H;�>�0m�2X�����]��\�/PF����w�j�\י�������ϙ��Ug0�%�����=Nn�k    IDAT�˃4��Y��"�Ł���@O=(��V��2�6�y�#&�Z�8j�J{�E$�M@x�T�6l8�� ���s�ϖ-�������Ã�T��Ô AB��s��E��e�cQ}��Z� ���S�����"��G��x�؋����	s0ؘ��%�t^�&E=��3�Y����&�-���=��*I����M�������E0�Q3L����zR���U�V�߸�	��d�q���UG�{��j��G�$c4���pu`y/��t�U@�r�dAXP4N�ε]`�w���l�W�tf�5�_�ڙE���c�g� Bd��PgQV��������������s���?��-�����"�����ܞ=ROO5�n���7�7!G,\�o"'3��놝�)5H2e2��a���9u4�3��!5 8�xVxq/��˼;��G��`�>\d���
�W����FA"{�f�jO��k45�hxh��>u�P��������G�Y�L�����APo0Z��9c���(/�e�갲R�h���9�&S�>���;�G�)�DBP�=p�	^���:�̤�}�M#A��z��.3β�j{�g���@}�x�xԩ9���I��a��=���l�H*��%: Z�>��o;]s�5��2(��� B�����3��DT8�44���^,V©N��"���y�Z�>
�gv�;���������I�#��R��''�a�2��k#�i����'=�������
��蘌^T&�H��*/=�N��n�R��SO͙�	��J��\���.��q=;�#����jw�N���-�>RhIN�uVݷ� AxpT
�1ֆ��p����k��f�ޣu@i���Z�:.ue�.��Da��brωr��Q��q��q��u1­�b�AX-���]���h�/�}��
^��"(:+��	�Ԗ������@��B����#N��lZ���S�X'�����@�5V�Z��г��5�yM^<"	S�i��#yP���0K��4��[���wY��XZ��KRJ$�v���C�$�[B������n�|����f�\��g�s�q�\Cs�[jw�"4����?�fAt���gW<iߘvqϬE&��<��('��Â4���"B�Y��#o�02Ȕ|.='�(��]5�I��J��n�E+Р�˿� �IK	E����!E���s]ų\�&�}Gu��q��|W�6��a���;��&�Wgk���=��C��S�B2����燫�U��+���t���SdZV`�l�O�}���$E;߯�SA�A!�gGi���f^��G�AEY]B�8���w�Z����6���;V���@����pҧ��ȭE=Iۍ��;d�1���	\�E
o������.��]_��ɾT���᯻x^��ԽO��@�1��<�n�����xĥ�D��k�ߴ6+���,���@�a�8��7�4Qf[��|~x�J�2���e �4�g��ѩ�]g[Z����K܅��C�A��W���'[�� \e��@��G��r?Ti��~�D�;[�ǆ�|�̻��	�!�L��m<���P,�ǈt⺪u�_t�D|�d�>���[M���@g`;�/U�:���6�zs������z�r#K���cq(���`p5jG[�
HJTS����b�z�$%��-4��6t��J�������#�m���
������B��5�C!��A���2-D�V	��/��߯q�0Wo7*"����?r�oi|��x0l�����v+g����gd�0�E5.�(�U�Y��6A�z���卣��pBq�[�eF4Q�Kv[Un�D8�;T �����,�X Ti!�#HZ�&,�K�<�u0J"���K�� c�v�!����y��!E��W�m��|5mA�𝌸Z]}ʺ*1~b Q��	�Sv�]�F%�Ҩ4���/�q ��R�8
��Al�M�#�7a���0�Ã�ɑ�>�+~���~�0�����������9���i�<dF|�)c��R���f����s��q���G$־�ݙD%!I�l�or�&b��i-9��D��?�{����I8]�����h�&�H?������ 4c��~��j`壬����+Yݴ��z�lL	8|�SLT��}�'���H��������9|V����鳯L�! ��{��������Mϡ`
*�e��V$8�O7�=�g=3W;���Q�M���3��o�R�,�>p�;�xS*��g�^�j�g?���ѹϰ�0�ik���O��p����]��f�V�ǃU��'sD���{�=����Ue�±���-�2{�^H��� ۆo[���m�����+�_��EAA^�U
�����!(ĿBӯF@^��?*��紉�P��:)��/�� ~����n���N����öQ�*�H�_F��}��!,���bw��Wۖy��}deQ��\C�`h��(���+���_l�N8w�Sد��E�6��%�6�e�§#���_K��R�v�O|��Or�?���7�-�a�*�z<GĹ |�BL3��D���c[��0�u��#�������!2��J�G{\\\GYY�ί�.�
T>}�lE�F�Iʷ?�M�N�o������$���ةA��E�f;��L)Y�O�a9�6}w�,��on#�\�P���;P���x�����/�u;O��ZC}�&�~�������;ym=YHZU@
��y���NOG���2: ���̴}�v�6��7���"d�(#���h�&Z0)�X�_��v|؄�N���|q0�T�P���A'`��0z_Sɻ�X���C�f�m�����
Y븀<��̠n���t%�	���d�A���)/ e
�US��������nMYz��v���Zf�D���s �*p܆�n��]�N��p<��� �����]�Y16�OpQ���.OIl�sM����п=7R����g�iv.�o����}b�gr��M����>��C�i�mq��6�: "�ɢM�jVH��,�}&�f�H��	U���q�]-���͉��70s8�%�dq�+ű�j�XY�x/��5m��;�����8���������?��B�ѝأ�yI����"�m�y�r{G{�?A��N��}��^3eR��"q�(t���?hP�U��a�&Q#3Ħ���E�nN�x��'v�&U�۬#W�Ϧ�\o�sa(�k�Gh�O�T�QWS2�Eb�zB��c#��$C/����(�v=v=9���u�Z1���G�Znj�G\�Yp΁��wT��U�H���:�#�BP̟����C�D�����u�׿v9���F��G�U x���HV���j\WM��a�-��G�I��Ԙ��-m��/m���UP0v�,z��>a^��Ⱦ�z?ز��S��e��Ci�ĜK�4p%]�N!�d�Ϩ�BW ��k�����(_�V3G܄)��5�Yj���!�b|"ѳ#���UTTދ1��r��2��kP��N�i޾�$�I��^�A좰�.rf��`��8i�*!0�y�?X|q��6�IɲV3��{��O�������y���x�Y%���=����FoZd?K�~��
�����C�����{A~+���5ӂRw�ٸ*�F�o4�7'�{ �{�N���Y����O�4D�^��c�y���"�Ju9%W��ra)��]2���z�!��D��Я0���<�x-�ݷ
�3zܐ|����Wh�x��\����D���J��AyEx�1@�(�q�c�1�C�[!V OK �C���*����P��И���z�� >.�ht��R���%^�@ no >LE%��d��wx��<�)N�y�04>®�|q..E�I*6`�����(�Z��^k����w:�Yج�o���KF��-���GP�X�uM�c����39@b�����=��� ~M��G3�l�?�
JX����"��5��ʡ�w�vC�&!�2��Yu�����wһ���j�ޥMoy�/�� O*J��ts�x^���(l�������k���.��������Z�ގ���M�%4�3�p�+����c����}��8�����µ������l�q����Y#�z�X�������T6��1S�������g^�u��j״�a�_i2�5&Ry b8�?���i���QLݡqn	D�/mZ&�3eS�zJ������;7�<x�N4�Bj�b�w����|
`�Y򐆈~�!T{�i��{��]D��.ɼɹ�zZ+���!�"aJfQ�}��/Gc�lAP����Fc��%���y�ڀ�����ii��l�7���SE��;T��Z��N��p_ޟC����x�hg���J��m٥�;�qr�R��e-%���xO�Y17"h\�F&����:�.yT�?���Я-�K�S��'�7��
 PQ����#�Ty�9���5PJ(� �TF�����F{p���x���M�[D37~�i&��'��Mrnʫ�v��B��7I��c�ޒ���_����j��j��F����}1�`�x�'�v8W>��j���2F�?
����
FR���h;bo3ڀ ���wjh�m@�yS��qV�k�;��2�m��1���W1�p�����7�����8�K�۴���&�O6�/��h�f�����<����}Np��N�yh���9~7
y�nM��.��K4�Cc��_F��Å;���(*m�^|�}���2��;A>Ç�,�t�a�s�WD�EB<�� $�(��^c2lyD��5�U�5��fW y���"�quޯ�+s<���A/W��֝��3ٔ�5���p��Ev�ߌ�^�TD�-&=��+%"�k..�Q{/��B�� .	���"��˰�D�һ5�W�1��Bbn��u���{X���rD��o$�t64I
�pV
5��ж���Ñb�
�_��'}�vd_��2��|<S�Bg��>�HV#���4�v"s2�g}�xu���Q�,;+�<5X����ż-2�* �jܒ�Xy�zff�v�v.B�>��3Z�}o{���*��8�z���eі��ڙ՗[��8�h��	@�@� ЙI]]�!�����A�g޽�c��#����#����z���VBՒ��]h�n��//��	>7�+(w6���ƣACcu$'=j��V0����&��'Q��)��"��6��0XP����D{��ǤrQ���QX��n��g����e�{%`?<+E�	������ID.+D�,d���պ�TF�^L~�^~�A��^�#�^=ZV�	O��pS�=j�DF���-�1X�H�I����#�W��PS1�����z��.��a�a]u�h�@���;i�.P�<Rx�>c�<rr���19EGu�l��X:Q�d���� ��'�Z��t�g��'1��?.T<��X�V��T&&�2�t����?W��kȬ܈�K�n�S�;y��>N�%��R�N�[�eL&�|�H�O���{�t�D�h��H��wyZ�6���T�)l8e�ǭ�v�ʂA|�&���Do@0�juʠhI�y}fja� G��a_@��^��Q�����M����E&}R��T��7�,L�pS����l�c}r+u�r�{�{�]�5������(.�&�ޯ�	�M`<f����A���Z����~{c�������	"'ᬳ}���67���L��g��ɋ�ɩ���%��Q֝�&;/��eb�m͎���ެ�WZ�5��?�7���|y����HFF ���>�Nm7μ�a�`z|GB�J��v��7�$3-�i�����m�4!�2��\�O��x� Aq�J�m��$ͻ"��+��f|'�u�
�6QH#j�r�QM>jV�m� �<f�b�w~.e�ёލ �j��*�5-.g�1��ss\:�3�+O�|����!L��K?�m��
��毉��׮1�q4_/�1
	�&���yN�,�%C�F#/b��;�b�`��X����I���֣���0SK�b6�p��a��0�8�/����w~��wL�y��5�Rgo��^^�(ѹ���:��I�[@��Ո�a�[�I�ZӨ������j*�|/��x�\�+׺^O�雏'���dф��ao�^� ��T۽%��An�������oS]�el���}����~9�s�f����!�F5t|x�RI��L�F��O%c(`��A�O��|:\ɸH���7�&�X�z5�R�di�$��>�6j�������s��A�$ه�J�{������1�<�N���O��2�J��Z�6u��񱝟׉�OA9��Z�����|��lط3S�(��ӲK�NMem�ƅG ���=�jX|�URr�r8�"�&K��\oU���XU�O!���u��(~p�PH�|V���T�s�ƚ?>����A�)w#����nԭ5����LW���z0�0�"�8{X!~35�����~"%��ӕZbU��.��3���eKC�Ro��/s�i��zA��j�]?�Z�� %eX&�b�
�֗�����8�6l��J��� %��R31a��֞�N���IT`��]��Ĭ�H��W�j�2�V���n�h+�.���7)�ғ!�3���4AT����&.�7��9����~�װ�Y��ʢ���ќ�Ƥ�B�,ee��@lWHj��mE�	��G��3�.���\��EG�'�w�o9-�0��s��{Z[��C�jh�w���K����S�>��an���3��o�o� �fW�^�	��d�V����R���<��P�C'S�߇B�lBV�p�� �:֗���V%or���mݥ9�]�h�y��2�G]qndBs��L�FO�p�G"*���5ǝ����M-��W�|S������\�'�u�BQ���t��8���pu���˽&S����q&5�v�����Y�]�'��Є�w�ʒ��l�L�Ge�S�����m ���[$�K1��X�Vu�ϖ�Q2�R�g�F�ކC�ّ���_> x�Y�p��ͽO����ș_���fLUhfH;V#I��[1�(���IM��˽��B���*��C����߄z�� 4D�葳���q��]G����z�;�'���.ݼ���ⰰ�HT ,M���`����O�f�V�寍h�6^A����(���t+2h�b
�"����_�!�h�JYx��W�ϵNyo�C�nu��>B,ۤ6,~;t`?���]����M@M]P���"x��ۯʏ�� t���T�o�P���3�����掟��0�1���tK�[�۶�Yr��D�~-B�&�T�%�u�k����l���IO�VA��6T��:H��	�?l�$x+Ov���e�S����g.Mt�3��K`ͥ��J�/�4�N��}0�{S��n�/��YR����� ��^���@��7y'��Q�T!��o���HU���3}A��d���y��K&�l�/��s�������5w@�[i���~�A��� ��,�3݄���	�6�f�M��ק�X<��m���~�~��X0J�{3�D�|� t��H�������)e����P��H?��O�$���g�>��o�oa��s���I���h��#��|��v�)1�,������;c~�Yj��}b�N���vK3��0�O[?��l,�v�T�|�sy�x���G"7�5)X�O��jf*W�y���ﭫ�.������t�Aliҭ+�&j)��1NB��((��=q=��nR�ɦI���2�rȲ��j&����I߸2gc	���������H�y4bY9�����(��w�˾�t��j���;�k�`dx+���{M�JT�������Z�l�t���|��t��\��&��}�i,w3]�c+��?l%���m�b���9g?%Yv������LV�Z�HϬ�^	d��������j�J��k��x]�E�n�X�E&6c������DRZ�i�B��S5���ug��Z��'h�NN�0����4$����\.�{ށb�i���h��
�Y�2��Wr6뎥$��M�0�7"Z��Rs4� ��Z���O�88%�ʫ:�����4� �g�g#-��ڎrӳܾn�Bax�iȷ����`H���ϓ��b��׷�7�J"+/0�O���N���AQ5j-�ž4��y��xQ	���$)��.�?�b<�2$�>a[g�s�����_��:���zZ+�8��g~k+�X!�*�_;��\������	�B/ �&��ө"���ZۂGנk�0��ڦ�_�KSM�`�>�n\�A$�mH��.�ؗO�C#.�AQ��Y��ZX��ug�<[;�ʴ+�?�Ow�x�O��VaH��u���⽈8 [觙�&F\JO��-�I��TӔ�[���E*�z��C @�	3K�>
�g��;AA�����\/�eԶt���F ���PmO�;�?�e�9A���o�ݣ��'rw�(�bA�֨<���Ű��	T���Tշ�sv"�x�UE��t�=�f\?N���KJ`�2�,5?���9������e)�7���P]�z��S���TAe{���>�{[�NYi��^�;8��D&��!���K���X�p_)����^��U|B��P�8�4��HڄT$��^�)<a]!A�7�QC6�������M�f���t�O	ib<�����?�6U���KѸ�t�k���`�%1+E3�`+1��+�d��xu���}��j���$�L��
lwH��IH�������5�=aݻYH�W� U���;�ꆾ�PE>%�*�hV��"L��L�K�!���3�}�C_��7]P�L�E����D4<+�Q��0�^yX�Un/��e@y͟o�B��V@���k�6�t��c�4�S�_� �!���(V�<��Mhh<s�!�t����$��6�L�¬34��$���!�'P�D��nm�Y�|׎h>��9��ƣ�Q	���5l�^͝˝n����*���M��s�y�Ț�<��JA���zKP"M�Mm���z�7��8�tA),@'S%ѕ��,*f�����^�����Xz�2�P�DT����.7(����e!X��ā����h��&S�����@m��Ra`����G4��	X�����썶p��[��ZQ�0�^G�l�E�����Xi6���Ե��a�"A�t!?���y���C�M��T2�]�6��"z��9�	xA��F��lq �Xx��X��2l�c�Hkƣ����5��3���.�J4��u�Z�����i�����]���e�`�*���A)/�@B;���H��9���9�L+�o�T�����B�f�^~W�I��M2��CZ�L� �U��E���dqM�&4	Ln=W`̮>/[鿜��2uqHQX��=����'�3����#WV���p��Q.���0�c����f�L׆�)ɗ�qv�70-ND����?_���oc�������+�D�5��'����V/��=�ً8��xy�=	ĿY�4S��Iω�ױ[�?��BY7�-�~6��n�lyv�Bc�pȹ�S�W=����t2	����hQ�0�S0�[U$�\���V+����Ի1�`��/�,y�y��,�.}b�ߴ��6e�@����%ˌ\n���,�~��a9ޙ]Ow�!�l1jN'}F6%ڿ�6�M��/��XU����Q��ʸ��\�8r�z݆�?Ӓ��R��k��3R�h>��'�N'�~26P���d�5�t���nL�uj�$g�q����0����E��]LȰjF�X��_dB�����K�w0�Q�(���/�m��y�uQ��V���M��Ѡ`-�1̏��/:��"c1n!K8�I��*�	5U�����l�L��w��x�u�Ug��v���VZQ]\'DgK�]���$�T܏��Zfh��U·�L�E���\����M,-�HӡtǱ��2c3O>�*5}t�SL0��'<s�hB���>H����%ѷ(�H�V�7l}n��XE<����~mx�n!�&��Nc��7����s�b]#_��m`���J�����(�{K�����6p�F����zv�������a������t�l�9�ǍͤUԺB�d��U��G@�s�h�6�����4� y��H��6��Iȓ}��ލMN�95��Qұ,\�]���fY�yA�������zB�I�b&v]k�=5�[�#,�^�(=IjjSd6��:�b�^S�RR����D	�~|��l�* ��!pB��h��9��A�ԗ���E{S��E�Y.lZj�H��-o;�8J� )��gL��$�8���D� ���X��o�?�?�����XL9�����'���Ŷ�S�5i��Ki?�b�ZʑV�Ϣ|�t�4N�<��z�|G�����'ex]&�V��C��#�t���;W1�a��֎�ݝg�/6�[O���}/�_�<
.�1�җ���H)P����i��-��t��Uf���t���.��9t�J������`8)X�i��F�џ����Ki��{�P<��o��@E�' B�H�k�|�?Fp�B�a!���鏟�1ǆ�{O����\�~��K��=E��B�AǑ��]Æ�=u9K��Ǵ�x�3�?y�3(�4�,��B��!H����H�I1�I����r���L��ڙh@��9�	�g�A!:ӱ�]E���"�����)FeTdZ`����d���xR:�\��me2��g�h/���^%�A�Vpu�"o���䉈�][4����X�l��ѕ7��qG�T�zd�$��|4="�wR6K��T.�c���&;�Y��xb��&*����ĸ��1:g>_O��K����?pg������'��:���x	�{���z��Ͻ䃎J,��\Ř�ңp�UL(v���j���7���$;[�/w1/�A3�lQx��������`%�<�/ey��C��_�� ���]r{�!ou���bM�%�Fx+�+��8�K�3�ML��S������h���c��?Ѭ�:�[�7�s�P��Bw�a�I���g������>c籋(tl��W��x�5�^��M����r2�Wm/ @�EU�-1��܂�r�ՐM}�v}9l�iB�P�1_^�ȥ�j�Z��+8�5�kW�5f���!����l�վ�ǃwZwY�eB���GH�%���A�#�<X�s~Os�s�E�Hf�!cL����l_8���
���ƒ.T�p̶����͹��UN�}�gߚy�&���%�F����Ұ^�Q@7̸�����u�X�Y����Ũ�y�T_�(R�TD���)u��t�!���	v�9��HZ\e����c[��>����uq��|(��iO!�R���8%�	[^���C�B&H��H/T��&[�/��Gmk�s��w}�N:�c����� �fIrZ͟�X��S�˫x��Fep��'�� ��r$�#��H���Lt�MI����r�ػ�l	���bl昳\�y�.��s��%��a�젾!�s^/�J�V�ݜoZ'
�;o�{��a�!(�MN��I�;J�u�X*$S��#�/BF-��t���˂��cg̽4�y�d����9F��2[_�N�j����c�ź��' �k�EN+:���v b΃��ƞ��,��C��䧺���bR)����]:��DV�2��<j�3+�}��V�/���.�)NpW�����y��G�|��kևю^���jj����"���!y��h&N�T�A��aL����Д��E�M��k�Q�	�ma���ȷ<Hm7ٛ��Oܨ�R��w`��D�yF��מU��X�2ig,5B���Rۓ:e���3p�װ�y	�TFC�otJ���D(Cu������`��6Ԩ6��w~Ϧ���\W{�IT�|�5$\�֜�x����%�l����3n�9]�B�/�[�au�����G��W28ԝ:P��􀲿��dv=	(Q]ˆ�̥�|;#ЛG�t-hw����"�,��ؗ���Y�!��(�+�Y�O/T��Td�c�����V|M�*^�Z�OcJSNo~i�'>��;T��;�ؿ<BF��j�@��.�1,�������l۫��2��w)k�jٿ����Mg�7VOX�)_R�p�<q*��۽��K�������:v�댍>�%)s{��8R����א�
��R㫕�Ɲ,��.��!��t$yfI��y�)�ϧd����H5� y�/��"pN2�z�jF�D�^,���;�G��#�|Z/��q�Y���U����8"���ЩA_E�Vʄ0I��ʡ��V!����c�h^��������9"�1�NS���Rʤ�Fqُ�� �����b'[T�W�)��ʢ_� Ӏ#)щ<�:G7 '|�����&�T)�G(c��nZ|�����w���g�o��T�6�~X##�3�A"�ԣ����%�W4�/���E4Zwa3*�� �T$I@)}s?��_��h�/y�(HߍOq���6V4����r}`m)v���$�j����f,�z��؟�ǲ�XYm�y�est�oLdq��%����x�˿!�Ϗ�h��E��ͣ�B11�&Fء�i��O�%��]����R3�
	�<T{�k���ȭ)Y���%�l!]�-|W�"p�{�AL,~��_�s�\~4���e����{��m��-#v�!����Y�!��{�(��|��&�� W�U�I�nZ�� ����;�������~#i�Mϵi��bfl�-o�>K?)���$�n+��䅴������X	��L���A���nޙ��Ɓ�i��N�X�mk�X<���+��v�;b���4����S��>�����=0��I��@H?K�D��#,,���T�TSe��m�[e:`HX9��E�<�K�@ĭ⅋O�[�FJF�Yp_!I���E���i}d
���qd ��MSD4c��<	eT\*�
<��qC(�I�6��(�R8Ii<�S���w�|8Hi}
sA�CF�|ü��j����_��ܣ��A,��]�O��*gJ_������b@N�5��1d�e�+���M����1/!��f���O8h�)�G�N�n4Θ��.^�tVԬ��C�p�~�>�b��ewK��mL^��Eﳆ�~̺W7��o��j�?� o�F�q�^Q�P)G�=��X.��<� ^C94�5:)�*g�s ������ Kx�X�e0��XH��!e�j4�߶퀐�����Z�ttt]3JfSi�+���V/?��tq���	[&��.6��:��_��o'��->�3	E����N�e�ϫ�S;O��ܕ�ʰ�K�|5�b���P3��rGB_���W�&���o�r$�\!��]���kF�&&�%�'2`��5j�4���E���à���K/di3-N!�'�i�nRaf�;��/���;p��}�����^SU.�6���:v"�p-p��%�I�x\g��Q���G-�eb.�M�Y�'q,���wj�Nb�9il���W����8�1�G�V��].�_��mSs���h~$��+����BS� ����٣���u��uY����@ $j�N����R� �c�\�ϙA3r�/Bv���(��p�d.~���l�Hd���*�?��l<\���?��:4�k��'�[�t
N�����!k�9�`��Bԋ�E�NZS��Z��
�Q��0ey��]�n�UQC]I��~�Y�:���Z�e+���G�z{��BA���x�%a-�����7�,�-{�����>�Sс����@.OQ���"�ߪ��GL�V��Q.X�6,H�E1:�,��?�]��n̔�R�SP �H%vˆ6��eF^����=��W�m��*{#�I�Xb��>�|ĭ����wa����ED�ȫu[\����*G�Gv%*mkΕ���O��z[9���h���tFHy]U�=#ַ�Zg���mVW2�A��Bر4�)��W�tUH =�:vGySd�d�8*� �bb;��;��]���!�6þN�m�D��U���T>�ƃu�	魖�.H)nF��)_�x6���3�
�ztu��vq�(�΅�Y��^Uf�g���o��L����5�����
�{6Y@0��WKc'�sE{�%�s�������� :d�]���P[ύ��\�R�M��-�Y�2	y�/u���D�Q�hW������_�J���bF{�]���>'\��5`���&9)Z�f:�?a����������5C��D��A`2��&������R+qki���/j	�b-��/R�\1�O��m1:����'\YH�>ݑH���͸x�K%��ȴN���pI�khW�Ib�O��"̺�E�_��kG�k�%�����Ô��b�Cz���1J�:z��3N�h��w�{��N.�̮��>%6���(�k��p�HK����ƜgR��gZ�x�)����(�fy��/������T,���e�Nm�|p�v��9Gz���DW;�T΃.R��	feNp�2��N�Mt��\�"���[�����X�"M���Z�BZD�pe�sm �"}�j]6���|�IJ8�:/��t2�ϝ@Ԁ���6�p��@��G[@x�b��FEO�����lo��ϒ(���ۖ�ޡ��զ�ºoNcޓSS���WW����wȧ���Q�F�����⨲���7�����̽꽗E|�bbyxsH��wZ��J���̐�(�O�ͼ����`��]�en#f'J[.v�l���XZ�4:u{Td�8%����ɪ-�-~������]�dLo���2�D���/�B�����E_c4n}b_�=�����,��mw�!�����D=Tob��kj�-�|�>�>j�c��M�d���^r7��b<K<�$���N�p>��3�|�6#� b՜��yጘ��oj��pu���'�DmP�)�<�|i_V<K� C��M�����-F75��3[AC7�%����L=��p��1~��s.4�۴��2��~�'�Jw�$���S��.��E���W�NJE�1L�=��l�x('j�FD�w2d�����`�]\�9��bAg�*z{.���JA�Y�%v�mk��-�w��J�ۚ4Ka�
��y�7���z��[��R_$�s�T]�.1�{��kKZ���{cq�r<�KC���(�.����A�F�`ơ`Q`�7�A�z�+g����H}Q�G��* t����6�R1��(8�~d��������@�@�$���B��q?��7Ñ+{#}�s��+� ��И/�7���������/8q��=Ƃp��u|�.�i����.���#��Z�f�9�@E>ȗ9Z��;W��	
�&Qx]@��΄���<�]�!��,X+{҃(eS+�l~?�y�1�rGEW݆^�??�@cLLP�0$"ҷ�?nrDML��H��e.�A���W!�%�	k������Oc	�x�B�u6���3��k��f�m~�[��'�9�",�x,�����v�q�.-��g�_�c��~��k�"��g�l�}�a����Nqh�x�g4Й@����v+�p���q2VJ����y�<�~�3��ѫ�pM+w�p�B��_^��Ā)WK����MI��I�>�"��⅛���׵$P�>�4*Bc���nL�̎�t�F3�6*@(��C���� ���䍞�|��7Ѳ�1ZԂ�[�_�B8�I%j��*�&���P?YT\��e�L�u�Ϫ��7+P|"�Y���W�v���zx+]�W)�h[�1��ܕ"�����(=��L%����y�ɀA]�OM8�	%q��b2�i)��
����8R���m�V�@=��z�:b��=�s����@lY�
�TR��<�K�`�����`�h6�]�	|Y��|�0�?�V��!
��$n��n{��P���4�㌐X4��R�o�*}WLT�>[�����ۤ����%5 �21�v7�;Y�k�f��@`�J�9�d�Ǆ.��|x����s�7�Z	J�t=fV��5b�;��(Fn��v�;g�@��0qݤ��Bd��;�M����|�c�O��֑� U�@�\,V�d��������A6�z��Q|�ڪN�(9�f�Im�Nk�j7�X�g��M����B�
��ڠ�"�7b��:��J�AB�{�=���ǉ�ݵq����c�$V/��J�pŇL�琖o���$C��s.
�ۨҩo6@�4����sY�Y�2�笭������.w�)��ꍦ@Jl�ݮT�M���ݣ�n��	b�p����t�nt���>��R���.n�U�� �l7�A��a�`I>Č�˻Cέ�2�n@�o�H
���|��Lk)�8Κ��"��}Mڬٵy�1�~�S7��{���\���w��������,4NM�_qm��^>_�U�Z�Y�X��l��~�d��tL_�iUW��w��U`9F�6�����qݨ�BaG��ғ��d�u�3�C����P�6��J�k j����ȓ�kg�����8,�Rx;� BG�������R���B�hm�nE| /���.��SSSN=$��_�b߹w�
~Y)�M�B�κ��ܨ��?/�O�S�s�oZ��AO���W�^#ܒU��3��:������G�fUQ�M\��,I�������-y���%���?�N-Tnj��7+7�T�7�\�v"d�ʊ
1f��v��uS,f��2�o�.;��͠`0L]2���+3����.�B����L��J>i,�U�����/dKA-�v�����B�I��
�1<�^S~��N��=�/à�#��N����O�\����Ь ��xb�܂�٥xP�{V������I��������SZI�g+n��1϶
kҠ�)q֙�]�p4��-Wf�o}ī!��WEs��֌sLE���L���2A�FD�ٿQ�O45���^�Q�L��i9� \Baޤ8uW��L�s�d��qNUS6�JiTgT�ܓ"sa-XTOˠj�L�@l1�VH��	)�W�ΦD۔�/�lu�U���i��"4���SB2})`y�Hl���Bc^V�<�cpJݩ�`���}� c��c˚��7�S�BI��"NU�G�\�VQ�E+��C��D�e%�qz	�^;[v�3��I�L�C�q�YHf��rQj�`���z?,���T$&�M^{���n����s���E���B�]e]��/��}i��\��[\����*kE���B�mcG>��D\.s�H�����P����u��q�mAܵ���)q����-պ�M�����q���TP�;���ʝ�;~���)1��)�%������3o�֐m��}����#wO�L��� �vT�~���		��? ���l'7�W��2 9f� �4[b�z���)%ԣ�{I)����� �@]��#������!�-���J��c�+�%:�m��f�(ez�ߜc�YвV+>���s�u�fn������I���Ul�P�)�ǋW��賰_�2L)ʵ��Q6�Ax���gw�	/���M���C�ݓz�L�S�'�x\r����×f�9�a �Q������FC"A�N�b{�=��M��`�_*�eD�[J�S��Ԁ�Vdg��9) �EG�C�ފ	w��eAF�a�I��!��� k��35c������D�k8՗	R��;�.��b�ڊ+rrl�Р�
	8?��g����x�@�)Bl�S�N8!�?Lѕ�0C�Ĺ>�KN<����x| �� �+^������g���6�M�Y��0Q�����we�Z�@�0�
�yӛޔ�w���纍���u��s�'�9�~���W�����`�����1xŊ<��L��9�Z�^~�Eu���r��}��Ҽ]O�/���ݕz�V�wݞC����Q�kH�@먭�FO+�� �#������/~q�n��D��Q�
XVҳo�]��Z]�r�E= zjq��1��@N+c�� `F�S�=u���q9��Zt�����O�Ld*uۉs%^�v��d���Tb�Mh�Ü�!q��Q ��m�C��0$Y�\88����~zf�_|q>�{�J����ʤ�Y& C?D&|��_����Ȁ� �q��B��b� k�<Ϣ�Qv: �C����_�>K�<����`�1�'�@�K�ӷD]�<�(�L�����!v�$ �Fθ%R��aׁ0Lx����h��=5�gR�#*=ݩ�ڗ�w[c�*��2r1mrT� ܞ�KePpב�ȱ��S#6#��T�
fZO�0�3U��t�i*���L	�Q*�ؐ�T��
�#3U�3�2��Vj�v�H;Lq��Id7|����wU��{�Ȅ�n�^�|�3�fˆ�@��9�����$�=Lլ�� ��3����͟�ɟd��������h7���p�'?��p L������
�I��rl���r��Z~ٯDCv\�HƫK�2+�`�H��"F�dR4���Mg��9ޕq|���s�,77���'<;�Bݩ��|ڴZ�.�#��~��[7ϫ��ݖ��&s[ޏ�]�)I�49NOdU�21�����kF[��h�TH%`d :�"L�LQ��Y�:���0�9��t<^GpSs�7�8E��c]�n�Yb�f�L�>��U9Ǻ�םj�Z�2�O��3�,��M ��h!.���`��:�b�s��p�3����&�L�Q�����.���Mٜ�s> eyZ�O$��K� E�J6:�@���;R�%��Y�83^)��Z:�xvC������F����\���rD; �9G6ie�����t�v�:0S%�6�{��QV���e���eW�C{b���vU���d:Ʈ.S��og:��:y\��V��} 2��ѣde�X�W�.d��	q;˽L��i��_@f��l<�3��,��9ޫl��g����8������Єa�0�hw6gu���~�j�e��z���-�	�@�=���.�&6�@]M�c��ϻ�p�C��e����jh�:�D��||+�����j�[��s��Ϧ�(�	�o���|*m�
ǲ4�5<���'\�����#9R*3ǃ�d�ѡ�wesmw}q�pDs�����ɮ��+����eH"�>��@x�W�Y�欎�������m7]�J�`ٲ�/?p4��4V�9 ���ifG�*owꠑ��iL+�a<m�	��ɴ��9����R�w�39��X���Fd����9��3�@����+��e�Ɠ�{v�Fv����b-����J���m��I9n,���~�}Fg,W�]����I�^$�)^�N/PD�HA�qz'���1����=��bW�^f��ٛiVciP�-_��h���>���y噒}(Cd��i[ATPҾs�/�jH��r�w�R�Rc9d����}#�R&%>�,6J;��V��?��q��LR��Y����O�]���p�#�n�|�p^���1'Ǉ��3�&G��:T՝V��S�q	�g����f�i�H�S��2�3�g��_�~��h�ZM�:y�v�S>��?���.�I�2�`�{3p�vY�q���t^�R��ؗ���<I��x	 �|Wէl<�|,K`��͑��s���f�`�mF0zw�R�̺u�N?��#o�H}��ʲF�	�� �մ��E��)�^RW���E��hd��v��Y�x�*�����r�:�SnU�~ou�V�G0j����X���#j�婴���-@Ff��;2j���Z�M��yO��+���X�0������3<�(�,ʤ�2�7��U�� (�-�c��s��n�|�p��ㅨ��2>��SfZ��y+�G�h�܋�1LE)BQ>j]�u�V�G���j��"�+�ɛx�`��f�
|Zw�f�<������FS����Rw*l��L���7��T�]�����D@x�:δ���f�QS��E�7c��]��}z���-���c�N�X����""A���N�v`�ʲ�x���׬YsZG��	/������/oo��;;��c��Z��<FR��]5`����`#����>d&��d!w���ޛ�Kz�����=�<d&$@�à>8]8W88!��H!�	(I��4�� �E�0	����9W�<xQ<�	��t����I{���ߪ��~�vU��ݝ&���~�v�7�o�w�����w����C������Nސ�{��4�?���u��Vq2Ĕ�|6i�B@��^����`x�&.;��>y/jy>c|v�t8�s�i�u�F(�Lޙ�Z-�z��R��J�Z�>z9���8.u��aWX��b��vw�*��6\)�B��w4h����� ����;A��ױ�;󌶣��+l?PF��ڽ�a[)+,�x��ږ7��E[�X��$>�P�U��;N���p0�r8�AaP�;��fo�?�~%��ˤG��L��a�e��!�JNpƮ�jc��_q�[�V�;kl��OW4f�&wD�I�v��A��{��M#�+<�Dt����r�2��xm��GOS�WG��6e1�[�v���	n�;��C����QX�������̵��8ײ���SO�N;�����9�t�DHT#��6��T��z����2�;�t�q�{sv7IPt�YZ��M؝��
2�����בN���j�2��x~l_;{���t�lo��{rڹ׋$"��*��vsH�bt���k��*�����Η, ��6]�f��ދ���G�T�h�����L�jc�����O���\����0{̭���?]�i��ARw��lg�n�j��޿�`��X5gn1CЬT��Y�u1�/�h�Le��.��iԢ"�Q>¸K+լJ����^�J+ѐ��k���wΑ��y� [��,��St)�n&�<qW�����ò�Z�m�W���w��q��2��`�إV3�F��|��<��z���w��P�o׎V;�z�Z���c���!��\/���{Q>�8�]��22m)��=��k,�m�Q)��k^[6(��l��`�,��F#񐱎���^�l�2�Qqb>�a���MY�{�s*�r�HHr�V��r�V�]w�UW�jI�����;n�̺R���Ä+�RzԣN�L���l��/N�H�#h��ei�y!8V���e�s��;BEG�!�d�ܨх�]D���&�.2i��\)�1�G�^�@X#��x}^܁,v>�5���#덁�����An�K��ۭ�y!�]/v�R�ee8?��^b;R'�(Ld��@��<Z,�'QI���c��K��!���ǳ �<ܯA OY��m㦗`��b<��B��s�$>�ed���G�х��R/r�~�oJB��ȑ)K�|^��B@z�AY�s��&c7��"P���|�dL�RO���Au�wl;S,�f�v��M���tZ�Z����v�EK�O|�N*m����q���\5=�'-_�2��-K�{�/��ǬLS�>���rG�0��Ep�x*������������.�hV&�����'S�Qʘ�a!4j�S��m�N��`#;���\��+�� l|�7x�r���y8G�F!����������EcLf�r��B d��c,ovfoԜ�VK�@-���mJ�F�tZ�Vj�j���p)M�v�n�<Q��R��g��ZKs�-&�Ʋ��q��Z8�>�ff�a�A�}�iD�����Bo�kE��s��%
Μ���
��[�Bd��3�+�[��a�ڼ�5�=)r�������zQ^��Pzp�n�Ȁ��00�%c�a7q��wq��{S�uAuKH�	q�l��v�Z�^��˖���8���K��u�KW������M˦V�5����^v^Zw���h�S�Ioy�1��L����l��	����IK47��7�^a� �ph��Բ��z��YfJ���Iৡ�%�G`���q�?��@б�.��>sv$��q� &�|@'Sj�H�����{$\���`��9���2�����K=��d�m���s�Lw�;��� ��	˝Tj�ScvO�4gR�4�j�N�R
L�?��� �K�T�J��e��)�jm�9m���|���Ԛ=�;�8;��@؝ǩG���DFL�b#�=�.��Z8�>�od@Sk�ހ�KP���~a�7����=�D� �;!G�9'�+j�(qu�m�p���ƿ��N23�گ�Z|�%���ʖ�CdO#�}�g��.qv;4�&�-�)i���C�R/�P���duR(�,�[R���sL��ˎ�o��S�{V��I�Ӻek��g�����J�l�9�l��
uD�*�
#����/�A��R1��#}�@�zq*�J�0HbM�9ݱ���0�0�s](#�I!H�����8g�w �IƉ:F��4�ܫ40�IM��Y2���:-�b��#��?FFbor7ctb��Ip���:w ѭ��)�k_��\>@��_�j.����G?C���g���x�X{ww��>�y�/��?.�����4���T�{_�vfS���Cw�T�ו��y�;�SO�e+Ҋuǥ�D-�|`w��W����1u=將����B;#O0���P�7o�^ �F]GF��ɹ��ljp�%���A�w !�ƽ��9�k�17d�K��#�a����e�l���	�-����}�k�@�?�����v��v�n:� y�k�naͤ�$g��@���7�Ŀ��/���u�s6Q8��s���ɓz����IEo��@��D��z{^d�⊍K�;�W]s\���t�=w�]۽s�Բ�43=��_{lz�K_�V�_���_�����D`o��N���@T���i���A�L�l�� [#_(�4�����Ї>��R�1cr�4�>�bg�,��Ʀ�0�j�AS��h?��?�wQ?$����<�0eư1@� &�8�@y ;�b||ϳ��]�ʝ1�5��n�������
x�	s`0�3���9i��N>�Բ�bq���-w(�g���Z�6U:�Ԝە��ܞ�voK��L�4S��wC�dT�Bڪ�Ruٚ����R�0��d�g����O~*�y`W�*2�4Y��obx��{k��`C�Y�\u�U���漋/���+z��&��n5m�?ڿǩ�9~W��N�y��6b ���������}�O�ց^!yzق�~*a�8��>�M��A�z����&������ۋ.�(��+��r>G��ӟ�}0��乭�a�T$_`�7���_n�Z�J�z���.wē6}��t�Mo^��g�n��2�RJ��~��t��ek'�?��?�;��Uw7j���ac&>ӹeY���\v� �mDu%�*�
�qC�#{>9":s��rC��h������p�0W\qE�����2'TР.���h����y?L���2���svW�%�<���tf�x���)����n�|��~���;5�~9p.4P��戈Nw���=3�3�} �ukW�jj�NcWz`�m����4Q��r{&����F�of~�rjWji�]MS�O�ם�Z��4ۮ�=Ӎt��@15�-1?�K��s�zPF�3	�ِ�v�=ٰ�}9��/�D�p�����'�5��0a�Jr��y�X����c�3F!p,&�7  �����D�6��3S.�4�ͩ��:����U^�n�����DٰU��5�\��i-���og��>���c�9����{�2�mL���� "ЋqǲpH#������2����\�iӦ��l�r�;�5۷���]_�K���w��?��w�ȳ�j#�QL���]-K��ŀ޳[* ��>8����7\$a��ѝT�<�Q�A��pܓ�`��@�k;� �E�t��(����.L�Q���t[-#�lE�ar��<��S~�2[�Ȅ�;����� � �lي4���W{�9g��kV�j��R}O�ǖ�س#MTfS��Y�n��@�E�Ze"��Ժ����N�ʊT��Ү���k?��y�� <37}X��y�`�.v�� a��QA����:�������b�N�	���{���\_�� ��7lؐI�2����� �eP@���r?���9���F-�S׀0�� I�B���b�S��(G?�����_y��z����#���1�K��u���;���hh��w�<�v��n�Q/������a I��z�D	ڕ#d�����O{��r�Q��S\��q ���(r�$�����1�"x9����սa�L��U]�a�}d�N6Poh�	:. Lgְ���k�M��e���.�4N�c� a��{Lx:��Yg>��{���r=U�3��Zy�-�$=f�e�<�f��ij�Ҳ�'�fuEy���    IDATjt���F�����;YK��Ls���ʏ��Ud�9����l)�0��Z���u��g��Äq�e�Ev���XU\G&s� �er�~�oܸ1�=y  �F��"���[^���~�ٸN�]���ס��s�6H�ֻ�޹�[����/2a۪�^O*�%c�yb���/]�}�KW���(G��Z�利5I&��G��x*]ȇ�� !t�8�{��g&,
tL��^���Jd�g� qɘ����?������KV��԰�);F9"2�x\����p ��f�6�=1^��	+G �c(�x�;�^O/�[��%�޶�0�VN�yu\^��`��3^�"���J��g���Ք��� �J�SOӭZ�\��4�^��Jiz�����S���v���j�?�m��� a�� �@8�罅N'�,�r0a^xA��7Оq��Q�X�r����BL8�����R�0����~{lSc�x���{�gF�H�����C�0���w���c�0��@��@x �B�:����K������ߗ��q!j��FG�h�DG4��R��b����3�<8��m�*��|����W������?��yGe��ʥ����p�x�2]EA�@@��	;"jx���"ƀ1@ga�(����a��Z9B&� g�#�ZV�a��.1&@8�NV�#�h�y�E�1=���rskV�j��R}Oڵ}Kj��@�5�Քʬ��p^�����J��=:5*+�\�H{�&|mᩱZJ�V�m�Lx���G;*���d���+�� ��V,[�`� ��0a����=�����*`L��Ӡ_�=��<[��1��g w�8�#���b	���w�0�G���g/{�U�~����9"t����w�ؖ[ߴn�֗���3��!G81�z��Q�T��dD��3q|<n�F�h;�c-ch	L�0�^A��R�V!��� LF��C�T�`b� ����
�v��d"�	kP��Y��݄	�LN��	+-��9�L��}r��4��)�w@���v=�K	
L�e�Tji�UK����?�µ�go�����/�tA���$���~X�/��E9"�	c�Q���)DQ��Z�N���	s���Q�9By��F�҄#����
��Ș`c>��h��-�&x�2?䜋a��r&}����Z�HȜq>K�;D���> �D�r�R�0P\)W>�q��Y2&�o�r��mY>��	+G�	�<����y�Atw�Q�o*
ed�a�0a�)uc~G��	#�S��-��&���l�P1hX/S;��&L��LX��r� ,�	�	�|E�ӯ�<� l]'�# ��R� ̵��N�9p�/f����l��gow��61��# �j���s��m����&<�A�&	O���=}�SKӭj�:�4��ѩQ]���X�=3�>�'�H�wޗ&�*Y
�kD�]�y8�� ��'抚0Lx!�s�	S�h�21�u��"fg����BrD$&��RL̙��? �L ���!!�� �=�	�Y&�g ��N���	D ۧ�=��Ȅa�BB��	wCtK)]�eo���x�8�kA
�_6]��v獗��~��k:��r�!j�	3� �0#��ZL� &���}o>o� ��R����f�a�R�Q�U2�Sa$�\ef��n4A���@g6�� �L�Ɖ��QR�����K�;1�=r�W���R��+>w��$%���e���_si_�/�gz&�zr�Yg�t�Ks�i�@��4^n�rk�|��	ۃ7Y� J�SK��JZ���4���ԮN�F��=����O\�vݿ3M�Є�~�8���]>+�	AXa��1���A�w���0�	h�Z�����W�l����8A/�&l�@(�/@� P�/�cC}�����%��`BX�K ��=��RF��sW�ƍxi��s�� a	~���.��%�n�d��7�}�D��Fs.k�G�X�k����w�9/֨כ$���>��E�;l���S:-yT8�'0�όV�D�<u����9Y�a@
��B Lc����]Ӹ����;\��o�9���c�+j�>����\ <#*�3�%��;�񎮜#t,+��,̆�}��O��O������"7�w�m}h��c��@0~<
���Q��� ��^���k�涛k�s�=���H�֯J�V+��{S��>�:�T���$=dI놪�"�Zf��jj��Ӳ��R�6����|`W�����������R�3.�E���6�J4�Ձ�� �ع瞛m���f}��`�=�~�d9̫@����*^��+%$J}q��r��r��/��x��!MG��^q�_��aꎸ}"���g��7�pU&�|@�Uϕlp���:+�5}vA}��_�܉I�&�ўMF_a�"��[��Vf�JLeT�奍��L��/a�s�  ��+קs�9{�����F��P4����T��K�g*�����6�����??�Ӏ�Z��!`иѭx�k�PG�<*�5T�����p���x��v��m�c��ѹ��+���3�����q�����3p�7#��z�wup�� v:	uI�v"�r�,�@�R�B6F@0�7��l厲wzw*wHu�L%�O�	JC���vzrn;uJ�t��.�)͗�?$�I�����gg�\�,'�!qζF����开ðW%7�L��Ja�Gam���{�mhk��[��`�\��z\�T�s�|��U��|����+Qh��Sڟsjȁs<��(a�+'�B���;/ u����_�k�\�?$��B&���	��sR2aޕ4)'�f����	� ����m��ǰ�{�	�G߻�es{s�	�	Q�'W��swo�'��< F�ȃ�E�Ӈ���z��X5B>�|�+�7C���Dy�T@9�YN�`�#�tw E����BY�{;���n���\~^4�c��5*#8�g��c�%ǚ��e�<��kG�<���,Nf������ێ欲J��;���r$L5�X�2Bml,��͜f2wn7G�3(3���R�CFo��vE�[#3[9uJݝ���rg�Tx^K��l6�� ����9��;_!�[��ڹgjF}�,g؏	��I�eb(	H��r�e���1#Iq�s햿%�c��R
�k�>��@�}�Q��s,�IP���2ǵMٵ�9��dE�"y�
���s� �sAl�ޭ�'l�믧�a���.�b�'\��u�-7_�n��,�OS��e*9���5��;�� L��
$8ډ�ج�4L-�M������H�{�~��,��Ÿ�[2p�<�09�k��w��ϡF仃�#�����������Ռ�P4b�se@�!2x�`Y)�@�=ޭ;����*j}�2c�Q����dڳg:w�����]�_��J�(l�����xNi鋏� 2���r7��lf<�̴�e��i�T��;k�ژ:q�|�w޵m����i[��AS�4�^+�B��-pm�%@�o%��mS����$]}'�<���8a>,�K�����9DGy c0c�/����"������[W^.��PO��sb��˲�񪫮���SNY���·�t��w���>}4 ܨ�Ҫ��U�ze�#����Dt ����o�v�cX�#G@�u�u�96f���e��m�y���hn��Q@ΑLY��y���)�=���4���"��Y3�]�0��s�G��2;hɠbB"�*0+KP&Yב	��b�֭�
p��1��m�x�,GĐ�ٺl�,h������>l�=�z�}25�����fNٓY��a�|􈔥�;�M�eE�q��H$M=M�\���i/�BU��{��s�;��2_�U�e��-Cq@�?���j>�y�s�9'�>Z,Rk� n����\�} ��O��&L}�f����,��d���F�	��c{u��+����3�8c�bLr������fn6�9N��/H��N���{`>D�Q0����o�[��u���+�뢱2�����?�gBۘ���'?9?)%��9%��&	���$`iL\�g�E���02Y��׭�ÌP�Qɂ��80(?Ȗ�`�r>��f"�y�^2�AL*{�;�ZwϹf���c��ɚ-�h���p� A&��[���;ώϦ�e,ԩw�F3U�D�/�AD�0�M5��Ko� -KS?��M��ڢ����� !����%l��%)1.��t۲ľ�v'�U��k��/���,- E�s=�(̗�)&�ɦ��+�����,�L�9��6�tؗ$�(��L�{�b�6�1�ܰa����~�]��<�>��n��<@xl�����E9�<�����֣̄͢��i�bG��#3f�W��ys`\(��a� /�1Ǣ;�-S�0a C��VrԈ���s-�@wD�����Fg��*���!���6��;��\��VR(x���a��L����>+�*���@�� �����x^|��k���|4��֟ݎ��N��8���gV��:�%2�l���}麉���C�8�AX�l��HF���CQB�]e�\_�I[��;��l#�g4�'��{�����ne�[��]I\��,_L�ﵰ}u�P�c| &���|en��}�c h��|�#�޽��� w�'�-��IY�񊃟�籜��Ah�!��,j`���6m�t�i��v�};��B˄�m�㼩ٽG��*�	31��lot���y�幹�A�҅���ő#dt�?��2aN cbε߄��b�fA��1�&�*�@�gu�ڭap2z��	|�}d��!:�g�3�\�<JCq-�����!"���xΑ�����!$�l�=J9�݂z�ϝ'�z�1 �;�ZBjH=�!�,���Y~�)�~�VsS�a�u�N��+��h��}ɬd�F���H��.��&���Q��DgP��^Ji��z�����w�C��r`'j���g��{>��ًz���JH�>��d��k0Q�¨�<�9��!I�I��)r�zDB �Ω���[Ǒ�Y/Vγ�l��ԽK z}������Y�����^��_OG=j]�7�R9O�,�D��+��y����	��0q'��s����x�.�O�8�1�]�����OF�ae��N����j]�!�ݒ����Ч���9�#��=�%�3�D�����' J�	|�A��'+f���$	��`@l19�9�9���A�_mI,9��7H�׿���9�����7.=fb9��LL�q�?�*S���Lx��`�x�1b��{dc���Y9�	��^3�?�����+0tm�;�Ły�\��
��`���l�N����?�:���8�4��Xc"��D��`�C��8̤��_�vԉq�s>E�2HT��IO.��M�6]��r��w�ly}�(V5�	���W��g�˫�ƪ�AX�(6Ha'�tK��t�8b�����o��[���ԣ���[����} �V"�l�8���t������9�> ��~�<�w8���m8������E���?��qz�1p�	J�?"&8�����b=쨕+'z�b���w5��u���Qwo{٪��Q$[�	��hPմs��4>9�(&ܯAc��j�`�:	e$��ް�aF+yn���5�����}�0.����}�5Qx�R���y��r�����#��?N��	n�6�M��~���\'���W�XLTw1�I�-�V�W*���#�m7�q��-/[��G��g"��j���6wg>��n�[���̣>�䟫���1��� Ց|�{�a�H��s��j����`<�����|�����]]w�u�j`��������Z���A��z� ,�ᤠ��N"F�̶U���,q����	L~�zr�W6n���%�# ᱻn|��{�z9 L�V�� a��L{oγ2,Ns�0o���9���+��V�P7f�~?21w ��=7�n��*�v�;��v�wys���q�r������a��;�j�+#�\�m$��(��|̓B�x������L���x���	��[��֗?�)O!��ȯ��,���nٚN�hw��Y.�(�u3`��[�,�s<�ai>Le�����1C�z��O�3�ar�~����(�@W&�pO���y�AL���_Gd�Ca(��X������g���ԐP%�w����3���?��������֋9�@��SO�:�^��A���ׯ�~��W6�fb�ݖ����Sg��[�D'�%,6�ofTn�+��=��w���T������[̳<���P��@\�{~̝�x���=����l���{��#g>���R�[c��,=Vف>�*��t{@9���k�S�ʠ�)�r��7o���SN9��Ŵ�� l��r�ZjV��)�R݅X��������X���`�����KZMFjK(���[��:���P9b1��	ˈ��b�q��A���\l{ŕ'��+5e���D�$�i�{e��_tԁ�ㇳ5��`��A�\��W]u�yK�y�ܭ7�~��0��c� �q9ڒ��\��s�6� P+��$��A&2�f�{8�ȽnE � �� .�D�E���8Y�jN@��f��u�����)��7z�#	��M�9��;�a�Z���j�Ì��uy��/���F{;��v�#W?R�k@Y��t��#K!y�@Ў��
eCsK�7y]ȯ�>+�Ҍ�in�w��E�nQ4*W� �,q$c���0&���,.۞�(��>�F;r�!�m\F���6B�g$i(Iؗ`����0�o������谍>�p��(���9���(�H]=L��+f�1<�p�d(��G�ɑXd�Er/��! ,�XH��VJF&`��y!σL8I ~�0s�-Yt�#Ev��8�r��0� L���y����g�0,@�\d8r��8�5Pd��0L��~��v�1�v�>$�1��c�̎7l��VaE���U#$GT*��]y�/;�.VZ�ճř�@�`�	;��	�9+G�	��Ȥ���!�mGnv��� v��y�a�h����!Z�u�
�醝.�$� \.��f���K'��	o}q�?���F.�/c �����_�żݒ��ѥ��@8.m�G@xXm��P�@�s���� �0a��[��;�dA�/���~�����!?��s!D��k��D$���	Ah��u2�c�ڞ-�ɺ��6&H���5��r-�0'�L>�;������ƖE�^
͌k��刻����hd�<�Y����[���y7�
[���.�L`�bbr:>�Ƚ�ޛ�u��s}��VH���7�t��`�����{mٲ%��|��e[,⹑����q9�^�B�R�~u�,Wsq^\��O/-ڰ+DM@C�L�+������ص[w�)�p�B�MxII{p��?�Wd��X��.}��gQ�I�e۴;OOH�LܐN�ܾ0lb����b�PW�@������'��S��T�KʱI�a�&'|����`"2CGgwדN:)�b�c���W i\�]��b�<��>��d�@��k�f��ʕu�����Ή���!7�i�������H?��?���_�%�n�S����1���V7vV�Ϡ�f����|�K_ʠ��I��^���];{�3��@�\}��Y]�'��C0����֑�� ����]��^�i�������`��D�;�=Ԍ�e�
<ĸ�2[���g�gyt�W~�~!GY�C4��5�{�����ڇ�T1H.��}�W.]�G�!��H؋���җ�4���+ۨX�	&�C�@0�������{���
�H^�WdVH0�w��]9��k���N.����Q��,u�cZ'q���԰��ߣ���i�π�Fa���.|Da�,z�=��[-]t�E�q�{\�A��g?���c����3��_�u����s];����w `�^�'���9>�{P=Yp��r�D�@�h���҃���U����3�*��    IDAT�SG�`��8�/x���J��|����y�>s�"~�gӞ�lL)�q�^{mցy.�����y��;+��>�����g�4�m��詍b��# ��L��Hq?1ȗ��e�	c��: )c �aN��3t�p�]�I'g��a\�}�{_ޠ�� ���
p�U���5_d'�Q��X�����2b:��Yf�Y뉎{��f��D�'�k�젋����~^��^l�~��s��l����[7$m
�������K��F�SIF��͠�WN�j� 4H
�*���U�
S��?�4ݿ��X����yW���-�{CD(�r �F��`�\�m�b���p ����R~Ҧ��Mw~�����������?l�#��&�@���8&�KÌ�&Ʀ~��adweS��i��?~�{ߛ�p��T+���<kT�AF�q��s���b���xc��S�_�T����Ox�2����:0&�*r Mg��;���5�I�y�c���|�A�B�zի2���������|%��;U3�������������ۜ�Q���m��sd�QۥLN��[���ҫp�,z9���l��MR�h������1�K�,~.GVjRb�l����� �̄'óAF�j$:T�;<�6X�s���W����W,Y*�G
cl�L춊����g�O̩
*���B.Ԑ�_�,2C#G������<�Ą@� c9�X��ʢ� LP�e��b�D���c���]6���>��Ol�
{O�e�����ԑ�鬀��/ǲ�9r������=���;rė���<ؙ��zg��nY��A��p�a�T�:�5~�9��b���.�E;�����W�-j�Q��3��('0/������� ����dFy��(q��w�v������o���F���Q����Q䚥�Q�5�K��W6o�|��S���!a 0�3�8#��I��[tCuU�����	�2h'D���p���ja\SƸ�b���9�=a�L���fi��놌�  �����0B��VO�s:$�#�L��(��ZL�!Gp�TF��L��q����7�1�9��������	�V��9ka�D��AH��`xb.���Aח�r6C�Q.��N�ˉ��ROFQl�Y�zV���v��6�F`�w$5'���<��z��ȤeД��2�G��2 ��W��%H���C���ny� &ܚ>*�SN���m���߶|_J��S���f�y�]u{����-:�����Ё1:.���ݗJ4��A� �@t��&�@e!@LGD{�����g�� a;���� ��_��E����#��֕n/�&���d�H	</� +tL)�����6˶�4�7�	�3�r���|�#�,_9F@�ikt�8�[���A�?���@�!��O��Osx���0&l=�~�!� ���w�3�atݵ�"ip��	�c�a< �w���k�ʹi��	��|>%�v!��y�(g|^�A�;v�P�n�t���Q��K���)���5�[~��uw�q����zXkֺ�����[��jz`)8����{;D�7�4���"�(�p7vh(�ݩ�;uA�c������9��>��W�V�	W4N h�����8"G�(���^���năB'�0l�PX�F�1�Q�_����!3e���o�g��2�
�<Ϫ���������8_�w�I��z-��;� ~��^7�o�+�№�ɵ,'�����p���?�=�FZ���N&qO��>\��MozӼ�<�~����0��'�����alOm�:����7d eҒ��|��w�ˋr	�9O���-]�G9�6R�,��^�[�@x�h��)�w&��pq0u��aus ���#��q��N?���s��<���5�0���� c�} ���+��vw�u��.�r�}[�w��9ǿ)|�����mGJ�ꕢ;�q�c-�Xi�� �����=��j[��O�
>$�����'Ot�aA�^zi>%^/>���x'a��a�D�7M�h�S_�E���l�)��wd�B�:���Y��:���y�[ޒc�9��,�S��L�B�����s$e������M���>��g�3E�0���z�	##`oN�E��{���afۺ�і� � l���7�Xwڅ �'��ڶ�@�����r�K6l��p�{��VP3���/@ ���Z� 
������eR^�cʽk�����0ꅻ��2acL
E��,�����)<��Q"S64M0��ו���F�TQ��������i�2>�z��B��MXu�yv4o@�mܓ�Q�P�����������/Lqnd�z%��Y���M������e�.��V�ݍ��H����as���� ?���̓�� C癉� zV����� �/|���$��~�_�'e��X�\��e�FNP��x�esPs.���Z{� �ddL�2X�p�R���.��g�qƶQ�b~pZ���7�{��;o�d�џ	G~�]u7��~S��v�0 �<ủu�
���S���;��;~�Cc 0����ig�`�w�V.g�3��Cc��I��θ�u	5Z�(�sm�=d�~��p�m�96���&<��3&���=�L�byY��=#X<qp����g?;����E&\�rw]ڊI?�vA\p�-b��vRʲ�@�2�6���^a�0er���9F�	����G>2ow��R^�-�ﬣX>b�#s�1�q��5»�6M��Q(�EmZ��kDy",�	�t� &���/��U����2[���Z��=����v76���Zٓ%`������J�c�k�ޣȾ�u�N9B}K@�5��0&�M&�p��H�x�f@6�������91��5�(7X�β���Ŏ;��
 Qޠ��� *���Y��9X������ d���� ��>�R��(j�N��J �����tz·5��Q���D��v2l�&����4��=�}r<���BR�;��@
�E[�ي \�+m�6d�!��'a���g2Yf�*F%$�E�*���]>A�ϯ��W�r�)�c3:�y�5�&o���AL��Z��
�$� ܝ�|�+�<R�I�n���N�Eᢻ!$���H:s���81' cp.���u�00\%��_��_�bp�Ӊ0NB{X�E�b[dg�9�Y�As�E����ɒ�D����Ʊ#PF�Mt������B������H g�yf�>�Iy�s�o� A>@X W"Xhb.��I�a�`;�vއ�b�+�㱄�!GD-1u��X�GT���g�-���@m�m�M� �d��0�'�m%4A��9ʤm���o��v�hH�� ��D�8����H���t��������HbJ������]�� |��/Y�c��與��0�l�{��[W.�N���I\;�n�t�ob�{nT�=N���ӊѐ�y_�E?�\Ɋs��jT�\�E1��b���#�.X�����ר{~��pbN�j��a�]��D�b���=��
��6�hA8ztN&�.����y���vz�Z�' #�������b]3P,�JF�MqON@��cT��n��X�e `b��퇁���֊ \�,�w�S����@��)}d697`���zaĸ����q1n��1@�xk0�f�&e�]B]����!%�9Qk���H�r���͛7_tꩧ�X��f a�3k�����ﾜ���D����{g_�Cݳ�a��h���}:�����j��0&�TV'��*q�Y+�K��K�cdE=�:���lK0�1.������jpAR�s��Nx�%�<(b�덢SzO���
/�0,�C��xQ�Pg��4`���d)��k��_	��Y��z�����;@�v
+���+%Y*�Y14[!��� ��N��z(��я~t�	��j���I�0:�y�hJJq��0�@38Q��-���9�F;pMV$���DB[uP���,�%�L��Gς�2QI&�G�&������}ǅ+�{�2������y��4��[*wR�\�����I�V'�:�<�Vnw�q�$/�
��o&�*�@�\�{��{3{zI�&�D��d�2���'�.ty&���ҁY�u�)�dŽeb1!T���E�w�f�����	1x�i�e�:7�M��1�î��w�Ȳ�w��璙��YR�ַ�53,~0p��0a��v�#�EpU�pr���dH䃞�`�nɵ-�sB����wK��e�,�!Ә��� �P����l��	�"���a�{���/�\�R`�N@�� �0���^i��IV�Q�ʈ��<�fFك�x,��wu�hoJ�@XFo"F3��\2�'�]�s%�+����磤R��H�zR |��͛/>� ,3E�貔V�}�4��\�䀵
����I�v)e�&�H�q����ie���S���Z����P��*ai�(�`? D�Ȅ� l�f9)#?��w�x#t���5��X���k6(uS!g��$�J���X���~@c2t�g@��{B�`5�ıL�8b�j�Q��<h��6m���O���~��3�p�,���gC�ޑ{��@�7,�{�"Pdi�8�� ��g���F����8�F#����q�!�D�VV�#��aA��A�:�^��#|�E��BC�U6
%�%�� j=b�Lގ�fc��v�-��ǹ�؆��͹A7����=~	G��:� |���ޣ҄�j�0�vW�7�r%�sY95a�N�u��*��\��.�J�J	�픺l���J�fbq��u=v���iPf�k�u��s�9#t}�������P�<��2��������s�=FP�ɢ�s d�5���\���ʬ�	�� �`����������5�&y�8�Ir<	'�;N��=����H;7:��td<��;qT��Ǆ����e��´1e�A�|G2(��y�����[z�ߜ'���Ǆa�k�x�`D�(��ނ^	�h�
!��KY��r�D�$G�������A4z�=Iw��2^c�9`�|ꌗsD�� ��R�t�[��֋O;���E�}A����[9�m˥��c ��Ċf .������ۨTS�\jͤ��z���U�ͥ���j��R�6ݪ��ک�.��c�fsY��^S�7V�z}��j-�t�Sc)��J�TM�TB�贲�� > &L�ct���/كF?�yR�mW1a ��LP��bd�fň`j$����0��)���f�ê�P�� �b�ѠF?� <��t�g�m�E���a����ׅ��ѝ�Y�����,��5�r{?����[zP���_?�L���y'�9�Aa���rϵy������d�9�LX��!���_�F?��p�~؛Ǒ!�&���'�<ϼ�&H��p�$h3�.H9鷐&���N�T�ߍz�9��c�)��ฟvUl�C��o�d��;фd�M�z3W�X*�����J�Ԭ�{R�wn|�����MscS7�'&��T���6Y�ٮ�ʹS�\i�&J�63	�+�����ޣ�ssO*��=��nWm��U���j��J\�ԕ'F�$��\Q���?��Og��I�/��8AӑV���NZE:SV���w��Y �(p��>�:�VC�]B�Ыђ18����Q:���֋L�2z�/���(.�1M�ɐ"���m�l{�e�꿾`�C�*G ���w�Ű��ʄ�7��A��0<@�d&LPCꢎ����Ya�c�鉆pBU ���٣��,�~ �@v@�brv�&̱ڇz���ԍ���^��� ��7e�c`�����AYf=���r�|ݦM�^��L��0��#R/��*����oj��Vj����3c�2�l�w[+W�C{j��Y>v��욙�������l���}�n��YY�L?��灧����(��i���q����J�N3�6�r��A�A �+�8�!Q���vt��F�㊑ZQ�R��+NRq:h42��������t��R>@�c�"tQ��%�<;�2�RM���#��Rl]�y츑!Z����o����έ{�K�ee~�{�s�m��@AX��>�iX��,�\x> ��:wlìuF�D&��h�L&DT�$S/z%�����`)��S3p��})�3� 9"�Dz�1W2�0�)e��[.p�D�µ�b��X�QZ�m|؁pK+u2�e�-�j�����Z}nrrkk���[��k�+�];��� C���sL{����v�|Nm��?9>��G&���ƚ�R�MN��#h�0#�E������w &��$KQ��;V�
V���t�4ѫe5�R��</�	a'k�+�RcVC�%)�𷱿$>gԃcdIԝ�9v��,���<����@A�瓝Y/� �?�`��	�3�fT���E&,k\���sBNonX�h�1�@�a����)<��A �|��^{2���h6���Ɣj"Qq��;X9��0�&��M&�aÆ�O?��{c/5��a]W�8Ƌ>8�e3��TN��DjW&��Junz�����U_k�\���cn��导c1�*{��k�֤��k;����};�;���g-k6�[֛�sqGδ������R'�zr�Y�Z��7y�n�����1���*�#'��D���iH-����$,� �� �l�D�;����Aȴq�H���Ag�I6�:`��"���@eaN�EmW�Q[t'רC:��2�������v�(�Y���eT{>P��� L����'?9�6��N�pϨa� ��aϩg!;�͌���0�{�8^ ؊9����Fn�G����w�oQ��;�x�T����<��?�	�Q[R~�;�xE���eMxes����!�{��H�r+5R3U:ci��2ͦ�{VL�6�f�[��]��1kn��4�5䨿�D�����{w\���Ϙ��[1^n�N��J�VjW:�A^��,���8��	'��9�4^��R����j"|�۷��]�y>�0��D��J���غ�46Q0�h���,�`���t,�����Дy�A��=�fmٸ�Z,���ۿ=����]��g"K^�u�c��.�o�狃���<��|�8���\�B�a'ƬdQ�����`W䦀չ��kz��e<�4 L�.��zأm�u�V�G\5�g=��*:��qo~繹 <L�o8X���L�)C���}j1vd��k&t�&��67�sD��y��{D���.���Oz7�����p���So�;kd�4�\��j��i��>�N�vܳ~�����zm�?��/ݷ�وv�c/{׉+v=�S�������?eyj./��R�B��f.�xg"��Ĺ��t��Ǥ��>+���X.�fi,����H��ܔ+C�m�p ��  �Ah&=hPFm&���=o GM���T��I8��2�  ��"WL��F6�� t�I����l���΋�శ}8~�7x�g�,����3~����j.֐-F���ڪ� `eY7;�,� 4�5�19�Xr�m�\k!���>��e��c��q/z<�����(�T@�6����C���84D��I�e�<���LDr�����3�YP��>t��҄#I`��J�r�[���2nV�	�ҷKS��9�5=��o�?z��\��l�����4��������{�}I��/XU�?�֜��߲�I��zf�0��]&�0��t�G>�'$��Ս�8S<�9�L_7FL�.�/��Ĝ�ј�)���?��?�,���.ai�u��0�0����1�W����y�%�X�Łf1 ���C���!Vv�le>G����$.3e�! ,� 
�w�w�k��q�@X ��q�#�u���X^m,�v;�G�_�d� h��I{��/}i�&��	pрIlO�RJ�@�X&'m��<��B��2�,޹���t:��箾���<�IOZ�dµ[���vl}���C�0 �3�U�i�9���c���=�c;O\����E����Sˡ    IDATuO���g�����w���ܞ�k�Vfó��J-䈉�x�� �1I���K�v�ַ��uV;L�C��#s�7�1\:�
�$�"�������&��w�+殺�̘.���1�����}�p�ا��� v"ʮ����-/E���^*-ulb�&7Dͽ8��"G�Ar,2.�9)�"��f��d &�ꫯ��a�N8�	�_��_���ш����)��@��E�������ZFuv�.e/ًԦH��	�n�5��3�]2�'M��wd�`�Oo��Qn=������yQ��7(?��uѫ�F�\���͛_��'?y�bl�@\�L�����̊�U?�����w\���`�}Ҧ.�=p�oMn�����=O��'+�v֨����X*�K���Ǆ3�k¬�۽����.ơE�"�L��;'2��8�AV����a59�.$@�}��&���4��t�a,8@�$�u��`i� 1LV�N�*;n�$�����8�?G�T�81����O|"���Q��y��8]H@N&� s�pm[$��l��F�j!9�p#R<&b�4��T\%���s6��jχ'lzMm�� �a˖�3\���Nˀ�4!�'�F���d��U������?�R���96�E�V�}vÆ�}�S�z�blv�&|�^�~���1�Fy.'`o��Sg�q[��{�Gw�]s���z�m�)����+�����tѲ���c͙��R'5K�y&�E��?=99rX01���5BfE	�2{�����(�N�ڀ8��!�Æ��"󛱔�� 7 Lg�%"���Bg��$t@����7��ܗe� :PM�_��A�p�a�׏�.F������u5�{���|�DD `$��%�6_a+L�E��k-���Uc�vŤ��7֕2	�c[\C@D��w�7`��`�b��=J@�rp<�g>����lX��; �@F��,V�Nd�>�&#k
v�R���ƍ_w0@����c�s�p�6-k�֝��{�9q��z���nԇ_����ZsԶ��M�}׹��{l<�K�k����m��]��DG�Kt�**y�vޝ��|��&�F,S�9Y���@c������ʯ�J�<�){n?�:2\-:.�K�q��=0a�4sNx�X��v���\��\�t'6��	�vu9�b��R��b���������mʅ��>`	p�l�� `NbE��u�Ġa�F^l<&l���@*d5Rx��a#8�	'�'�&�]�;֏�� ��&�0���MS%�]=�kRâ#�?�  a����Rٖ��x>=Fۓ��n)R�0O�� ���/��u��~����Q��<uPm�+��Єg˕�_w����?;}�	��c�E���n1�{�M�NW�?�����w��̩V}Y�4����I���p��/��3���cn�@;;�Fvg09����d"֗s\ygG� l���ς�7,�侔A���PF:2�� V��z���5!G o8��/�����l����\������&lG��]����8]��O����*1ۈv��`��9`'��� ���Rmu���(��?+:�Sb$�ep���\ĳ�l�76�A�9S 4���3�F��`�7eP�Xj�� LY�YڌVN{��K6��L� ��\�n���l�0 ����]�nH����������2&x�
~�����۷^\�v�]�G�*�6S��]B]��4ӣN~T:��3�X���������ǚ�UG$؁U`$]ѭd('��e�'ٶ�`�%F���L��c�9	;����G�e�^G��xc7���J�e�Pf��06�}(�0H��8���a5�خ�\�Q�})�sr�:������N��8qE�Xǃ���; �$��cӡ�Wd
0�:� ��[̑A,9�n�),�KԌ��
���@Oe�����2p��;@��q��s�OAI��I�H�-A]����b�Z�qP�+��"gt��w��kq t,u��9�6p^E�W�s�R�37n|��1�Em���,�0�]�Zz`�q�O���n���_��Qz��9eӻ3q����ݵ�7�7gO�V�v��*�+�Jn�N:!��ſ��kci|l,5���j]]�����t؅Ҁ�vtB�	��N��g=+O�D�Mfg��}��N':�M]�T����ݡ�/���� 	�����$���;`QtD���#�-Ĳ�E���ܶ�2�DPv T�z?�C���	{ �� Y�20��F���E�=�A���u�Yy~ ;�z���xGdA�{l���2O��J̮I�)�ڪ��种aĬ�ע���I�r��B���Dw�(��+��Ю%/��mذ!/��_�lk��#y5�����O�9�x~�՚+�˟ްa�	�2L���X{��G�~n����o�C/�1������;Ϛ����V4�>�Rn�Z�.�M*�N'<��.��rs�T���z��#� ]���^0�=s�J��b3�Z��h)c��#G��e�E0.���_��.�!��+�`5,��ED��H�9l���ʈu�`HLb�"u��bp�]�]��n���^d\��@�+S�z!����ds�>�%�� f�2<!@�A�$P֫�>mړ6 �hK ���Cޠ]yw�Rcܱ=mM�<���x��F}p.�b����N,bC������g	��\��B
EG80�\�_~�<�>T2���y�	K�[�"��������=�3��=v�-��z�Rt��^�ɿ���[~k��[^����G�*�Z�=�J���d��M��	?rb:󬗤j��*$���f��r���KC���e��x���
`�A0J�2�	�+�As�	{� ���ɒ��눎�B�saU�J�ɽ`($����` �a��2E�Ƚ�Xb�/A��8�q�g�}��f�e8�m�Cu|�m H�h�<�̗�$܊�>�'[Vo'��m@���H7���w���Æ�x9�c[��@�bsM��͔���[@S2��|HD�@d��v�_<��7�$F9����IN��v��="�a�0w���;8�=�u.x+ō'��6dY%6�;�$�	\�1?�i��A�l�����+����@��91��y�c>=��Qn~��YhZ��'m�n����dٖ[/[37}R�2Smw�R���*>�7�H'������Zᩉ��nv'��v{>�A����LBi �u�d�z����,�
�-��he��	�z)�b�iuDϧ̰6�Z����T��6��(L�g��`��ι��cȖ�*?;�3�I��I��2���D�������$D� ~�^�=Wtw�`�\�kB,���"�]��U� );k ¬zd�מ�� °W��6x&�Źh�xI��sh�N'��=�kڦ*�I6԰9VJπ��EM�kEF���xuf�}��x�����xhw�8�����ڰa��L����}B��{����ǟt��xMw�C�z�5�Ԧo�q֪-��Κ�=?2V�)Ä�U�J*��S���ؓ�����Y�@�hu��;�C`��>2R*�	;Y�F+@�M\�'� G���9�s�F�� ���r��������\�9@�8Sadh��f�j{ ;��E|%�q}&��0�v�������E�+ھ��n`<�yœ�~aꌥ耰��;yw�F�$t��/�b �=�7���t�#���jK@��L�~͹N��,�/�2^刮u���|~���}D	�ߌv��&.�G�C�6�]{��0����b���mګ�Vh��W��a�]��kN�������M������~����7^ݲ����l�t���*ө1¥4Y���N>!�uΙ�����R��������D�B�U��#��QtⅲEw����7���_W>>׏�8~.��,�w9�spY��5�% LP?���� "�ᚬ,lqy�g&FW�]3"��@,��Eh�H*`����3��������, ��F$�����6n�-Ѿ�%>Äq�ѓiC�Y��xC�O.�0LM�g6O�A����,���n=em���>���q��'��O��T�2�~:L�L�v*��se����(Ca��1�uw�y����1�R3�aQkV�s����kl��c����~�c7������<���󸍟Z9���WOn���k�{���S�5��6Wf��&'��U�צg��ϤR��N:�Ĵlr*���lwC��H\��]��6�52B�#)�����t�x|�C�]+v��Y��;:'1���V�	���9�������6��� 9�DB����;�%>�%�ΚG�x8�0ug�u��8�s���۫V��N�2t�Q�G �� L�	_�"�ri�G�6�d�6�@�k��6��b�y��QF3�2������a���Mm�gs���c]x��z��uE�NC������hO��>�ܴS`��!����3����}n~��z	����ʭ7\�~��W�g�n���I����\J�j����c�g��������L%v};���n|��m[ߘ��e�S�z*7fR���J�R����������/����Dj�Y���E�*�a��
��#D�#��{a�t
2_ѱ�p�C/�r�O�C+Pv▉��;�0 Ё	Q�3"W�v��vG}��g�	����/oT�ڟ�^�sd[2E�ⲛ �v�	�c�|T�Q2�����I `r��	S ��O7��m3@��e���@ȵ����=��1��,,bGp�+��8pM�E��j�� '�%(�;.tr��fH@,>��y�������D!�C�0�h�K����
��6�'3E�"`�\�Z���_�t!jh�v\��	��@��Z�j�S�J�LuC��?:}Բ����,j��RT�3����*w�������dgv�T�����Tnv�7�6t���T�=�ݗ&''�o�Ư�����nTD���F�F��AX�(~�;'P����P���x̀����
H=D���Pnf�)�g���Â���0/_��R�C&���D��sd& <�	kqp;��;��j���y3���] 󐛁�u��~ G/	ǐw���c�##�g,�׊R��b�ݐ[�I��3���(_p'yv�KYB�r�w�Q;v~������}�h�E�1��z���Qtnq�2��ā��Bl���~Ll�T�@c�Z�N��Ax�ƍo\��7^�v��� <3τ��~�<��Ԗ��<��/׏>������~ ��s�����o��_��{ǅ�=;�9Ѯ�f=3aB�J�Z��ȧ\M��qg�Uӹ瞝�y�O�Nj�z�;����1�+���;��E ׵uFZ�HqcqAa����袟;� �Ɓ�c�0��U�ݠ'�iGaY���+��޸V8���; ���s�L��zǮ���A��G$t!2aT�`��?�Êڃ	S�)F�X�~�b�c9�,�XO��9�- ��}�ss��f��}��)�xM����jM��R� ��sb��A��#�0@�����e���}����"��������9�������3E���6����M�ް� <vˍ��ٶ��T�M�R+U��t�R%͕ʩ^kͭ\�O�cOx���1_��Mu����~��'/�}�'w�󋝙ݏK�4�棭z��]�N%�����t˖�R�\J/;���'��͹41�l> �  ��y��0�;@d�<"F�v�^d]	�h���^l'�W�2�8����K�,aP>�r�atb\�Q�4T���L���Cd�����!0���EX.@';Q��B˄s��b_���= as���xG ƞG�Y�����߂�e3l,��`ɮ/l �m�`	pAg��F�oT�+%6Wͩ�82Yȹ6�AqQ�����0��*):!�)N�.��/��{�֕OH4�8@��AC? ��c��{�ڻ�]�����N���V7�D�r'uj���Z��}ԉ�j�#�����q)*e�56m*�X{�s��|�-�����R�������ިݚaX0Ӫc���'�����87����f�����w�`x��4��|\DA��ȋ���p#iB�<���X`Gh Lg�?/u��ϻ��������bd�0�1�c��t5����3 �V8F�c�Ja�_�n��P��.�l@���o��
�r8����w�3��Q^�+�6��K|,@(�.L>��m�u5_�-F���W�qxs�.G(��<�9y��*�%�u�,�n/��A�Xy��+&�)3 N���R�0\l3 c�\����p@Y���i�Ub%�_�u��z��z?�L�+�n����۶]��5}T�<�zk�E���DoM�ԩ�ӞT�4W���1'�oj��?��i�൜�X�cN����s�+�����s{�����i�*��ޖ�r�������4��ؖ���ү��/�S~�������T��r�8p=�d#b"K�E�sa$�0l#f����0��lh��ha4*߹-����u�`	�8@P$J]�w���N�ŉ�~Unǖ���Z'/�R�	��9�C��d��T^B0���vڼy���/ �<Y�-��}�M�CzDX1vc��h�zbf5�q��=����a�������zl[%.]Xo��)#�xõ���ye����9 ��C<��;����q�xe�{��>Pd���6�&�LD䏃L|�Ŵ��F/�߽�D�����eC@��0�,�T� �ϲ;o�t����hͮ�g2��[ޭ���RJ�R'ͥj�WW�gc�1�8��{Ձmq?�2����o�8�z�֋V��E+ZӵJ��ʬSn��'���c���.u���8:�Fz�ǥ��n��f����Ra!�(3���� \ԋl@����߲#����1)��VL�=��8 j�"���� � �	#IP&�W4�Q@�q�Ƽ����c*up>L���fۑ������(�Q-h�HGqr�g��mڴ)�2���d¸� :� ��&�8��.S.z'�_��O�m�Uk~�{�.n��GD Ҵ#�y�l��[d�܇Հ���p��v��l`㑈p=nX���_"�������m�6('�}'!x,���(C�] s*�͛7�aɶ7z���;jj��oZ����Z՘>�S�)Gnj�rj |��4��33�������cW���\p�(F��c�������<�����wl��W5�{��TO9�|��:�	�%n/U���N'M��R�>�M��jtݤ6�]@Ɛ^��e����Fo'���0V/��wq�.v נ/��	�zq��� �!U�%h�<#:�0&A�c�dγ��I
�B��Aw�ו>��;���#�At.�lLP���>�腗���W�` ������h��!u�{n� ����Ł3���A5�Y�0n��,�d�X~���|t%\tã�CS�y��(\5ʻ�2�z0�D&\x�eH 1"����A62*Sv���>�<�F��\�h=t~��>pRe�7��s��Ww�M��Z�]�r�L��f��j*�}|���Tk;��]�͹G�'�=��;^��~^w]�7l��t�g�߽������_&K�&�i�!�d�x�>�l��Ff�,��Ɲ�q��1�9�>�H�+��ҹ�4�� �я�c�, �L�bXLܙ~���\����OC;�w�S�I�{�b�5v�CY���Z�r �&��:z4����;c�A�:�SP� laYx&HD֓��^H�_�3:VoF�6����w�!^#�Ɂ*��L�+tRz��XV �]H��9Q��F��
�Q��Y�{�6{�a���8���$[��/���x�ٜ��� N��%�����_���-7�κ�;^��5s<q©=;�0aA�=�J�r�-�Ӯ��={V��������>��k[�,����������2q����w�󧦧?ٜ��`���"W(;� ��w��<Jw�	�J7�%��l1�Wt��_�A0C��E�l)�1׈/��|3^��b����͡;6;	D�0 �s�j.�'���)2�����s2��[1Z�/����f��p2v�A���k�J�  �IDATtQ�!u����"��4�5f{��V�c�@l�5��kjkʆ 0�a둡GV�5�������`��s,:=K��đW /�d��=)c������%K����ౝ��^���m/\՜9�]�M�v=U�K��.WR�Y��N���s�D��k�jc����������f�66$�tC��M�R@v�"�&2J?ը��q*hq��GU�6?Z	!T�(M?�&�*�
��T�U�4���!�/0^���̽��9羳g��ݵw�����̽�|��9�y��u�4SH�^���]s���6�۾Y��\ɩ���_o럟8�.^xP�_��?����u��8���BKA �q�тf,;+��t�@|Ǫc$a�lȓDH�C1P� �������Z�� L�<���!#)��]k�׆.=�	�9b�G�y��#w ������Z�C��]�����[�TSDK��-��3��N	���#�7���I��[�:�A�.��~��F>(����o+�F~DŭF_�lJ ��?�j�C���<=|5�Cz�vp���P�����B	=8�SY��5�[3I��v���g���?�	�<cn��+[��=����:ώ6ϸ��P3Ƚ��6�`:����,��@��\ԛ�zN��ު���,����G�vKc�TV����f�>M\z�M|tW�^�� �c��u����C&)؂k
�v&o	[��XNF`R@��gu@�5�_��MGd���I�A���݈ &�x�� �6M� ���@���D-4R6�H4C�Ǯ~�^��	�A�a4B��$)�r4�$��E��o�k*�@G�^}�U����y�\k �A�W� �)@���I/�2�w�JI��m��,=P� o�7�s�<2r#�����>�.�G|	���0ʄ'���pA;F:=�oS��	!&�'���?ڷo��o�Z��Ov杧�?����3�^e�Yd����M�1%{�g�����3�gU�����~�7��w�wYe�_�rx6)�LM�p��or����1�llL�f���]��ӫ��z��LN�U����hvz4Lj�%�0$,��L'��T�I��'�� `��I���#�`R3I�؊��.�`�F�du�����#�L2�0|a����(Y��?���э�ɠh��&�FPG���b��cF9�� -� �>�`���/�0��� ��$y�-�݂W���n�s��'�A;��yi�`�A:a���6����3�`��Z�.�v�$�?��0<S���;T���qz9vA�3 c3�%�K�w-���������_�+��:K�0��d�G�qݹs��W����\$y�z`��;	$O�m�Hpɐ�A&��ix��sΦ�d�R)�a��
�t}���I9<���=�K1d����?���ĮQ��j�M�PZ�F�R�ګ5ZĪjU��Ԫ��R�����V5�ؔ�����γ�z�s�3]��p��i��L�0�zo�y)@TYfvf��LS"-zDm�0z�EJ�Ę�y0P^�3�����=s�C["	��sPD8#���ﾶ�|B�����o��'	w��
�	.�S�<r�qҟ!��&�Rf?i��	��\�Y�N�mO�	$v��ģ�bHj���qE�ʉX�T�($E~���8�kq��~��s��~��VǈQY0�<��wm�3n�*e(��!2Xp)W(^FYȏ�M���ڐ0z��(���1%��Zp�À&�N�[���U�rZ��1�Y-E����X�:�%����Aio��ޘc&��g�����w?Ek��8�-�6[����j�1����?6ٞjW+E��M��q�F�I�6���F2�����D�< ��D?��������+)��n8E�	*�������V�m*����2/��}���$Q�� �+!���6h�I�5?E,�qI�Ʊ�6�:e���� Ì䠀u.n(=�f.oZ�*��ڌ��tZ�O��.x�*uS�ʩdKҔx+��$��ðc����:�ԸK�,��M� \����5(��k����wh�l��h�m��"�Κ-�Sڱ/�G�,{}!����;�~���T]��q��\���o�X!rB�:A~AǮ�w�ґ~k�D�"%ᭉl�4Ց[�<����3�XGP���:��[<��|^�8;�0�&g�7�K��8��B�w�n���aEߝey>�o4��v��%��4D�e�~Ʊ��?Ӿ�CM�5y��w�k�3�����d��%�G�o�=d�;���I��<�G N���v��<������0n�S����'� j���"�C~�Ñϓ(�<�+m�z���{@I���pY��9�qʇ
�#��O|n!�}�T"[��*yy�Z3�g�f�
����<��>�!Y�CF�����&Gk�sX�yy-®����2vW?-�ʁ����g���,x/F0��H��"Ax�Qu�����?�R-��p[�<���1�\�Քۡn�G�f�d�%���{�𞙅aF i��qee��#7� ��3��׏7���;$��iX�z}:��`�����LuB��?���<��("���y_���[9��ED��\�P��Q_!H���I���B-���M�B3jf�={�F,�7j�I�6	)�8�_V����>[����wkZiͨ+D3#�0��0���o��?��y�Ʃ7����?�?�:�>_��~�����Wn�J$����-�y�w-�U�!7�=�K���62���U�f��7	���	��I|���*,-�\eF�I�G��Q��x�銃� ���}�tW�B�� я�<�.s�վԣZ0y;�pE1��±G]�x~�s��duF1�T7�N\P�����K*�d�5H5��{���៏�d'O>���͎���xr�&�{�կ�B�;]Iwȷ�*{���Nŭ? Ѧ�Y�6���5Ɩ���Z�g�n�M���d��������̈́�+���]�&Fܣ3��ȝ����\��m�����J%�7�N.V^���lOI�W`��Ԛ�;��rFM�hO��&kSkwK�F�d*�=���e�yU�2J�~��s�<�<�m$�ȁb��A����F�1$�JCzG�9�0�X��=@��L\j��nl�˓�7��d��4�̈́���=E@���Y�����Y_ވ�o��N?�vҖ#b	�
�{�� %�R�o�l��u�i3����7�( �0_#G����W:�z�F�I�Sh�_���Ĵ-k	y�E����uh|�wrn�I���K]���+ԥU)�~��J�M��h:��,���0XyO0a��W�m����m�	i[p��������b�w,wk�n�i���2���|Q�aӿcOd�����ޟܟaP[_�BV!�,��
���I��ʠ�5W� �>���O1*��T��C�".C��±�$��&�^�o,k���`>������b�=`"���r�ʼ�"���T����n��րj�����B�������!�������Ѧ���C����I�ǯ���>ZHc�K�V��
�;	�`"���X
���/�����$�Ďv,�[��5�8��f!�-F�[i^�G��b�#�ۣBb?B�/_ɋݭК�Gb��xI�ݩ+��@0Z0c��]X�)��"����lps�lU֩ʑV
�&,��焾��;�E��sx�g�k���=���qH��/z	B�=���@�!7l���������Y��K��WCNC]�����:�0�w��0����ɻ	�%�e�4��()��c��+iY��l!{8� �j���%�&�Z0��ә�<���Pf��36?�[�z0�M�?���x~[�੓I[*�" ���.�$z��Y��f!1����>�g���D��UgΔ��2%z_�ֹ�\
���82�~Mg�kTZo�%s1�ˑ������ݣNw-��)k1��o�Z�F&WК����D���i�5j��W���r�mEwm;�u�`��IP����P㕗~��Ka����B0�A�q&�>B.���0בTI4K�� �i�?�R��1u�03<ԏX�7�˂%'�mj�9h���^����ivJ��A�P�4R�m^���P�MݸY��� 	3�ܩ��^	���E1�5� ��$q��lJ�O_&64��%*�����b���G��O�w��;�����F8P��cfpBiN�-1R<0#-p"ϲ���R��,���a�F��IO�sd���e3����I�F�]&�N��74}$x{L��*۸9��ԃsNVق>����{6�k�9�2���[չ��y�0�H�e�UKGd�V�)��
�?�R�:���l���<XIZ����l�j����A�h���r�W��y�8�X�;��쎈~�)S�v�O!��ێ}. �B���t&�Y��)zG�A�2y�Ÿ�3y�`�
��PeuW��.�id�sĻ���r������!?j�6�#ي�V��}�;�v��#7� �eqe=��q-MgDbc�,����<�=��]79r˫2���x3�ȧP=���}���u#AQ+��|��CQ}�Qűq�E���Ȳ� V.Y`�F4���w��o��{@���x>��	t�@h��;KmO+K�ҷR+��6,.��+2c��A����-r	��Y�����WZ,c�����2�*���1ۤJp�����h�J�������Z@�8�/ILM�����W�#�'�����J�|����q��ٱtǀ���Ϸ9��wW�wB�B�lk?%���������Κ�ꨭ5 �_R�F��Ԯ}�3�"��'?�2�S�t���(>����Ν�O��\��p2Z����4h~{{��8Z>��#@�Πu�Π�S0�.���sF	Pԭ��d��H��=��PX��x�v��o9q���="�J��[P����{ǭ����;o���NՄ�6��.��mE�������Ҩ(���<�պ�?	~�W�-e-6.�$���ɋFaZZ���?Ǜ������cU���!r��鐵�����ʗ;^';0i9fI���i=XI��ɝ���:��^�\�n�{7��>Ԋk�����>�;��Z_���0�7(penHV�3�Sx:�Ҹo�<��{@A�4�t,r�A���hqb�&�au=��S��
��.��E!��;\�(l
R�Tݖ�V�^�h����Qt{J�~aulM1��Z�'�}��:��~ϝz���I��`�ϊ<O�.��GS�؜��i���{�k��	�;�j���\�Դڹ�,`��>}M�=;?֘����D�bZ��"��V�aH=��ov��,w�pn�ө�o�Q�+�/?$U䴐�^��g�:ںf�c�j��д^�w'2�_�&.F�m8�z=E�T��|�����^�*`���r��.H|):�F0�ޟ��_�2���2B;���P�D�	��3�'y̭]]CGmIR�����B�|v^�=�}	�߯��5��M}�XI���n���2�S��ToO����ޖ��_E����KPɸ����Im���ˊp���D�l�"G�,cC_���G���)��ui|ۯ�u4�Q@N��)j��3�7zœu
���hPۋ������|�q-#&�1E�vK��/j�ET
#���A멃�,*-^�!��GA��T*u�*��+�6�6PŁ���\e4�Ҕd���x益�������m��Bj"�7.��̗m71�!��U����;<��o�]�K˰�u������������񏯣�S��FB��tC�_WW/鳇Z_� Ps��k�Ѝ��x �����ö�nv@9��s.ƒ�d�������%��V�C"��Y��n�qX�6�G�?��n���$>�z�c��,� �WF�.��}1�{����
W�+g�VK�Kb��6����w:Z�%�Ko\(�[�s���������2��=��($T���.q��hB�@3%��]d��a~~GIɿ$�Y����������k�*�[?Ceg�3��rƔ2��v���ގTڵ`�M�oOl��PK   Ȳ�Xݤ���  �  /   images/b275462b-1e1e-4e27-bbb2-300eaf3790a5.png��s���b``���p	b``�```��`�����HqxD30ĸ�0��gG�fOǐ�9o��w���m�x_��IY���I�'�н+�h={I�w���Kj~�������O��{�ֹ~��\�k�{����ϟܳ��;��v�{���wڹ�_f�!�=�vǼ�s�u?_f�^i�~�ߚ���W_�Q��lfr����ϓ���_W�|��Ϗ��?�& ݍ�h��{��땩����u24�Uǭ:�1�M�̯Wv<����u�����u����t�w�Ai�����ӯ[W�3�����k>���U�i����~+5��ӷ��@��vB�������O.{���ι'�����Ys=���>�
�.؉��v2v�5���x~�><q�ɶ�[R�乛��>�Y[XD�;�m���_o������mL/��ׇ�^1���{����Ǟo?)S͜������O*kc�8���_^\$�e���<Q
����}����U�غz���wA7��=:�-]�'#+���!�
C9Č�ǫ�װ30��9010t�A4����l}�������a`�!���� ���yv��ݯ�Kb*q&+?y����J��
$�Ǔ iB�\~>�'wS�3|x�������fw���Y;�
i�c)��\�F��'�v�F�r�{ν���y����n�;�{����g?r�Lg^l����+���A�]�xK����2���YZuUn]��Ҩ��ֽ�c�����o��o�g�6ojK+/))Q�)
�_�:�&���1���-%��OU(�~�85?�M��z�������;�+Obw���PGN������sO�����]{�1��o������+�e��͈�<���ywA^��������a��o����?���>����a�5���l�����{�y�d�ol�d�O����a&9��~.�� PK   �|�X䮃�  �3     jsons/user_defined.json�Y�n۸����ipH���ml�I6�Ţ(H�j���^�jQ��َ��D����ɖ�sF�9�3ҏ����O��ҕ�R��K���WW.�y��1YV�>u9<���ÏKs__{U-��j���G�Ĭ��y����j5�8Z�O��'��-�h���a�g$V.%�sF"p�p�)%\f�N��S�L�|��D�?~�'�;rN�,NI�c���k"K�$2�`"�Ƌ�3^�ȋ�"�O~��~�/3��l>û�q$ �x�������/>�2��d�*�+�8OoVe�蘲���2���g5&�1���1���ɗ�E�e^��ÓUYaRfƺ�<4��W�j����Q;t��X��L=CÚ4��L^兟��Yz��-���
�nJ�[^b���C�|��U�-�m�/7!�ro��~Q��W3�ֵ}{##q�NP�����_�j[~_���g���.�����engnw�tW�֋\g�Gm�*3ɪ*]�(����6�I�+V�� ӓ'�b#F�I��f��DZK��ˈP���Jé��&y��= "ݛ���u�����>%&��֫}��^q��^q��^q��^q��^q��^��zŻ��`+��+��E�^����smC���ۆ.&*F2E�n�1U�жA�,���D�b8�X��
a�ˀ��a,�h�����7�X���p��1~tw縻���1�_1�:���n:��+D�<%xߣK�����E|�?Aן>x	D� �������?�P/�j ��	x�&������a�~�5�!JnPD~���� 1O'�O�T3 ��D�)���=�(?ES�p��O�MM����%]�+��ij���W��"��k܋��g"M,#R8C��Q��}��Ԃ�G/�V�g����nef��Δ���j^�9��Ƽ6,���2!8�d;��itJeh��8q\������c S��#)K!Չ̈́P�MɃ�n�����W�+��ej����n�r~��Zz���|����/Y���Uf�)\0f	8p�c���Xu8�9�q���wUTk��Xf����55���WW�t0���n'R{s��I��,L���*:�0��H5�c�b�5"�2.���c������B�����p�&1��ށ҄e����7��x��->�ܤ�c�����!Oo�^�G�f�m���?��.��eۡC ����Ҵk;x�w�M������M��������i�v+�K��v�2����ܵ�W��=f���B�>\t��.Ն��t���'�G}!��cj�w�Z�7��?��[{�P�M:�=Cp��\�����Mki����	�(�d�Zo�o��g-�-8&�DI"HQI��dT� 
ݡ5/7k�����	�#<8��[ӡ��k�p���ԦD%Ѓ ��<6�/��dN�2KО9�R��=�荥�,�T�*y0j��Q���[<+�$��v��%�f�M(�� w���h�~��|��8.��9FP@�|�1��X~��8�>���������>B���׳×�� �^�g����?)lq=;�8���mϜ�u`�o;�[|�G����W���<��*�|����(�@��>��T ��ջ$\C`�_,�x�GQ �mC��A2LY�3�R2�`��N��}z����7�,{���ʏ����w�7�,{��w�vid)-��ߍX��Y������1����(k�bv��0td�e���7��b-�~����R�CÊ�n7�e���(��Yl�w�O��#��[�p��.��_�=�����?PK
   �|�X�`���
  �q                   cirkitFile.jsonPK
   �|�XG�~��  � /             $  images/0739a1b1-a163-452a-a325-ab452d55b136.pngPK
   �|�X��g  n  /             ��  images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK
   {�X ���s� �� /             ��  images/305f7d3b-a649-4bb0-9743-3edf8bc04acb.pngPK
   �|�X�B'�  �  /             o� images/39b1e261-4cc5-4406-9e56-f0681178eaba.pngPK
   �|�XhT���� ċ /             [� images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK
   �|�X�t� -* /             .r images/7a134b18-aa7a-4645-8200-8100c2fd668b.pngPK
   Ʋ�Xld^M    /             )� images/8a38ea7c-aa1a-4e70-97e2-d2d1d9cbf557.pngPK
   �|�X�Ƚ׌  �  /             Í images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.pngPK
   {�X��"�IY eY /             �� images/a366fc27-e5ed-4ac3-9d3c-a6e1ff305d7c.pngPK
   Ȳ�Xݤ���  �  /             2� images/b275462b-1e1e-4e27-bbb2-300eaf3790a5.pngPK
   �|�X䮃�  �3               A� jsons/user_defined.jsonPK      $  ��   